magic
tech scmos
timestamp 1428712110
<< pwell >>
rect -105 43 92 65
<< nwell >>
rect -71 25 -53 36
rect -107 -48 88 -4
<< polysilicon >>
rect -26 57 31 59
rect -96 49 -94 51
rect -75 49 -73 51
rect -53 49 -51 53
rect -36 49 -34 51
rect -26 49 -24 57
rect -22 53 21 55
rect -22 49 -20 53
rect -18 49 -16 51
rect -1 49 1 51
rect 8 49 10 51
rect 19 49 21 53
rect 29 49 31 57
rect 39 57 79 59
rect 39 49 41 57
rect 43 53 67 55
rect 43 49 45 53
rect 54 49 56 51
rect 65 49 67 53
rect 77 49 79 57
rect -96 -11 -94 43
rect -75 5 -73 43
rect -53 38 -51 43
rect -63 36 -51 38
rect -63 33 -61 36
rect -63 26 -61 29
rect -36 11 -34 43
rect -75 3 -62 5
rect -96 -25 -94 -15
rect -64 -19 -62 3
rect -64 -25 -62 -23
rect -36 -25 -34 7
rect -26 -25 -24 43
rect -22 -25 -20 43
rect -18 -5 -16 43
rect -1 2 1 43
rect 8 -4 10 43
rect 19 37 21 43
rect 29 41 31 43
rect 39 41 41 43
rect 29 39 41 41
rect 43 37 45 43
rect 19 35 45 37
rect 40 34 44 35
rect 54 -3 56 43
rect -18 -7 8 -5
rect -18 -25 -16 -7
rect -1 -25 1 -15
rect 8 -25 10 -8
rect 19 -19 45 -17
rect 19 -25 21 -19
rect 29 -23 41 -21
rect 29 -25 31 -23
rect 39 -25 41 -23
rect 43 -25 45 -19
rect 54 -25 56 -7
rect 65 -25 67 43
rect 77 41 79 43
rect 77 -25 79 -16
rect -96 -33 -94 -31
rect -64 -33 -62 -31
rect -36 -33 -34 -31
rect -26 -39 -24 -31
rect -22 -35 -20 -31
rect -18 -33 -16 -31
rect -1 -33 1 -31
rect 8 -33 10 -31
rect 19 -35 21 -31
rect -22 -37 21 -35
rect 29 -39 31 -31
rect -26 -41 31 -39
rect 39 -39 41 -31
rect 43 -35 45 -31
rect 54 -33 56 -31
rect 65 -35 67 -31
rect 43 -37 67 -35
rect 77 -39 79 -31
rect 39 -41 79 -39
<< ndiffusion >>
rect -105 48 -96 49
rect -105 44 -102 48
rect -98 44 -96 48
rect -105 43 -96 44
rect -94 48 -86 49
rect -94 44 -92 48
rect -88 44 -86 48
rect -94 43 -86 44
rect -83 48 -75 49
rect -83 44 -81 48
rect -77 44 -75 48
rect -83 43 -75 44
rect -73 48 -65 49
rect -73 44 -71 48
rect -67 44 -65 48
rect -73 43 -65 44
rect -62 48 -53 49
rect -62 44 -59 48
rect -55 44 -53 48
rect -62 43 -53 44
rect -51 48 -36 49
rect -51 44 -42 48
rect -38 44 -36 48
rect -51 43 -36 44
rect -34 48 -26 49
rect -34 44 -32 48
rect -28 44 -26 48
rect -34 43 -26 44
rect -24 43 -22 49
rect -20 43 -18 49
rect -16 48 -1 49
rect -16 44 -11 48
rect -7 44 -1 48
rect -16 43 -1 44
rect 1 48 8 49
rect 1 44 2 48
rect 6 44 8 48
rect 1 43 8 44
rect 10 48 19 49
rect 10 44 12 48
rect 16 44 19 48
rect 10 43 19 44
rect 21 48 29 49
rect 21 44 23 48
rect 27 44 29 48
rect 21 43 29 44
rect 31 48 39 49
rect 31 44 33 48
rect 37 44 39 48
rect 31 43 39 44
rect 41 43 43 49
rect 45 48 54 49
rect 45 44 47 48
rect 51 44 54 48
rect 45 43 54 44
rect 56 48 65 49
rect 56 44 58 48
rect 62 44 65 48
rect 56 43 65 44
rect 67 48 77 49
rect 67 44 69 48
rect 73 44 77 48
rect 67 43 77 44
rect 79 48 88 49
rect 79 44 82 48
rect 86 44 88 48
rect 79 43 88 44
<< pdiffusion >>
rect -65 29 -63 33
rect -61 29 -59 33
rect -105 -26 -96 -25
rect -105 -30 -102 -26
rect -98 -30 -96 -26
rect -105 -31 -96 -30
rect -94 -26 -86 -25
rect -94 -30 -92 -26
rect -88 -30 -86 -26
rect -94 -31 -86 -30
rect -76 -26 -64 -25
rect -76 -30 -72 -26
rect -68 -30 -64 -26
rect -76 -31 -64 -30
rect -62 -26 -54 -25
rect -62 -30 -60 -26
rect -56 -30 -54 -26
rect -62 -31 -54 -30
rect -45 -26 -36 -25
rect -45 -30 -42 -26
rect -38 -30 -36 -26
rect -45 -31 -36 -30
rect -34 -26 -26 -25
rect -34 -30 -32 -26
rect -28 -30 -26 -26
rect -34 -31 -26 -30
rect -24 -31 -22 -25
rect -20 -31 -18 -25
rect -16 -26 -1 -25
rect -16 -30 -11 -26
rect -7 -30 -1 -26
rect -16 -31 -1 -30
rect 1 -26 8 -25
rect 1 -30 2 -26
rect 6 -30 8 -26
rect 1 -31 8 -30
rect 10 -26 19 -25
rect 10 -30 12 -26
rect 16 -30 19 -26
rect 10 -31 19 -30
rect 21 -26 29 -25
rect 21 -30 23 -26
rect 27 -30 29 -26
rect 21 -31 29 -30
rect 31 -26 39 -25
rect 31 -30 33 -26
rect 37 -30 39 -26
rect 31 -31 39 -30
rect 41 -31 43 -25
rect 45 -26 54 -25
rect 45 -30 47 -26
rect 51 -30 54 -26
rect 45 -31 54 -30
rect 56 -26 65 -25
rect 56 -30 58 -26
rect 62 -30 65 -26
rect 56 -31 65 -30
rect 67 -26 77 -25
rect 67 -31 70 -26
rect 74 -31 77 -26
rect 79 -26 88 -25
rect 79 -30 82 -26
rect 86 -30 88 -26
rect 79 -31 88 -30
<< metal1 >>
rect 6 75 19 79
rect 12 65 16 75
rect -107 61 -50 65
rect -38 61 97 65
rect -92 48 -88 61
rect -71 48 -67 61
rect -102 40 -98 44
rect -81 37 -77 44
rect -59 33 -55 44
rect -69 11 -65 29
rect -59 19 -55 29
rect -49 27 -45 57
rect -32 48 -28 61
rect 12 48 16 61
rect 33 48 37 61
rect 69 48 73 61
rect -42 40 -38 44
rect -11 41 -7 44
rect 2 41 6 44
rect 23 41 27 44
rect 2 37 27 41
rect 47 39 51 44
rect 58 40 62 44
rect 82 40 86 44
rect 58 36 86 40
rect -29 30 40 34
rect -49 23 58 27
rect -59 15 -30 19
rect -107 7 -38 11
rect -34 7 97 11
rect -46 -3 -32 1
rect 3 -1 39 3
rect 3 -2 5 -1
rect -107 -7 -102 -3
rect -1 -7 3 -2
rect 47 -4 52 -3
rect -87 -11 3 -7
rect 12 -7 52 -4
rect 56 -7 97 -3
rect 12 -8 48 -7
rect -93 -15 -83 -11
rect 3 -15 51 -11
rect -102 -26 -98 -22
rect -72 -26 -68 -19
rect -60 -23 -50 -19
rect -42 -26 -38 -22
rect -28 -23 -11 -19
rect -11 -26 -7 -23
rect 2 -23 27 -19
rect 2 -26 6 -23
rect 23 -26 27 -23
rect 47 -26 51 -15
rect 58 -22 86 -18
rect 58 -26 62 -22
rect 82 -26 86 -22
rect -92 -44 -88 -30
rect -60 -44 -56 -30
rect -32 -44 -28 -30
rect 12 -44 16 -30
rect 33 -44 37 -30
rect 70 -44 74 -30
rect -107 -48 -7 -44
rect 5 -48 88 -44
<< metal2 >>
rect -102 -3 -98 36
rect -81 22 -77 33
rect -81 18 -68 22
rect -102 -18 -98 -7
rect -72 -15 -68 18
rect -72 -57 -68 -19
rect -50 -19 -46 -3
rect -42 -18 -38 36
rect -33 34 -29 71
rect -32 -19 -28 -3
rect -22 -56 -18 71
rect -11 -19 -7 37
rect -1 -15 3 -11
rect 30 -52 34 69
rect 47 3 51 35
rect 58 27 62 71
rect 43 -1 51 3
<< ntransistor >>
rect -96 43 -94 49
rect -75 43 -73 49
rect -53 43 -51 49
rect -36 43 -34 49
rect -26 43 -24 49
rect -22 43 -20 49
rect -18 43 -16 49
rect -1 43 1 49
rect 8 43 10 49
rect 19 43 21 49
rect 29 43 31 49
rect 39 43 41 49
rect 43 43 45 49
rect 54 43 56 49
rect 65 43 67 49
rect 77 43 79 49
<< ptransistor >>
rect -63 29 -61 33
rect -96 -31 -94 -25
rect -64 -31 -62 -25
rect -36 -31 -34 -25
rect -26 -31 -24 -25
rect -22 -31 -20 -25
rect -18 -31 -16 -25
rect -1 -31 1 -25
rect 8 -31 10 -25
rect 19 -31 21 -25
rect 29 -31 31 -25
rect 39 -31 41 -25
rect 43 -31 45 -25
rect 54 -31 56 -25
rect 65 -31 67 -25
rect 77 -31 79 -25
<< polycontact >>
rect -53 53 -49 57
rect -30 15 -26 19
rect -38 7 -34 11
rect -97 -15 -93 -11
rect -64 -23 -60 -19
rect -1 -2 3 2
rect 40 30 44 34
rect 8 -8 12 -4
rect 52 -7 56 -3
rect -1 -15 3 -11
<< ndcontact >>
rect -102 44 -98 48
rect -92 44 -88 48
rect -81 44 -77 48
rect -71 44 -67 48
rect -59 44 -55 48
rect -42 44 -38 48
rect -32 44 -28 48
rect -11 44 -7 48
rect 2 44 6 48
rect 12 44 16 48
rect 23 44 27 48
rect 33 44 37 48
rect 47 44 51 48
rect 58 44 62 48
rect 69 44 73 48
rect 82 44 86 48
<< pdcontact >>
rect -69 29 -65 33
rect -59 29 -55 33
rect -102 -30 -98 -26
rect -92 -30 -88 -26
rect -72 -30 -68 -26
rect -60 -30 -56 -26
rect -42 -30 -38 -26
rect -32 -30 -28 -26
rect -11 -30 -7 -26
rect 2 -30 6 -26
rect 12 -30 16 -26
rect 23 -30 27 -26
rect 33 -30 37 -26
rect 47 -30 51 -26
rect 58 -30 62 -26
rect 70 -30 74 -26
rect 82 -30 86 -26
<< m2contact >>
rect -102 36 -98 40
rect -81 33 -77 37
rect -42 36 -38 40
rect -11 37 -7 41
rect 47 35 51 39
rect -33 30 -29 34
rect 58 23 62 27
rect -50 -3 -46 1
rect -32 -3 -28 1
rect 39 -1 43 3
rect -102 -7 -98 -3
rect -102 -22 -98 -18
rect -72 -19 -68 -15
rect -50 -23 -46 -19
rect -42 -22 -38 -18
rect -32 -23 -28 -19
rect -11 -23 -7 -19
<< psubstratepcontact >>
rect -50 61 -38 65
<< nsubstratencontact >>
rect -7 -48 5 -44
<< labels >>
rlabel metal2 -33 71 -29 71 5 B
rlabel metal2 30 69 34 69 5 fromShift
rlabel metal2 58 71 62 71 1 A
rlabel metal1 96 7 96 11 7 Add
rlabel metal1 96 -7 96 -3 7 C
rlabel metal2 -72 -57 -68 -57 1 Z
rlabel metal1 -107 61 -107 65 1 Gnd
rlabel metal1 -107 -48 -107 -44 1 Vdd
rlabel metal1 -107 -7 -107 -3 3 x
<< end >>
