magic
tech scmos
timestamp 1427500770
<< pwell >>
rect -56 56 -39 81
rect -75 6 -39 23
<< nwell >>
rect -70 40 -60 71
rect -70 29 -47 40
<< polysilicon >>
rect -62 74 -39 76
rect -62 68 -60 74
rect -73 66 -69 68
rect -65 66 -60 68
rect -58 66 -49 68
rect -45 66 -43 68
rect -58 60 -56 66
rect -41 60 -39 74
rect -73 58 -69 60
rect -65 58 -56 60
rect -51 58 -49 60
rect -45 58 -39 60
rect -73 52 -71 58
rect -73 50 -43 52
rect -70 38 -60 40
rect -70 10 -68 38
rect -62 36 -60 38
rect -54 36 -52 40
rect -62 25 -60 32
rect -54 29 -52 32
rect -54 27 -44 29
rect -62 23 -52 25
rect -62 16 -60 18
rect -54 16 -52 23
rect -62 8 -60 12
rect -54 10 -52 12
rect -46 8 -44 27
rect -62 6 -44 8
<< ndiffusion >>
rect -49 68 -45 69
rect -49 65 -45 66
rect -49 60 -45 61
rect -49 57 -45 58
rect -63 12 -62 16
rect -60 12 -59 16
rect -55 12 -54 16
rect -52 12 -51 16
<< pdiffusion >>
rect -69 68 -65 69
rect -69 65 -65 66
rect -69 60 -65 61
rect -69 57 -65 58
rect -63 32 -62 36
rect -60 32 -59 36
rect -55 32 -54 36
rect -52 32 -51 36
<< metal1 >>
rect -69 73 -65 77
rect -49 73 -45 77
rect -72 61 -69 65
rect -65 61 -64 65
rect -50 61 -49 65
rect -69 49 -65 53
rect -49 49 -45 53
rect -59 36 -55 37
rect -71 32 -67 36
rect -47 32 -43 36
rect -59 31 -55 32
rect -59 16 -55 17
rect -71 12 -67 16
rect -47 12 -43 16
<< metal2 >>
rect -65 77 -49 81
rect -65 61 -64 65
rect -60 61 -54 65
rect -50 61 -49 65
rect -70 45 -69 49
rect -65 45 -49 49
rect -59 41 -55 45
rect -75 16 -71 32
rect -59 21 -55 27
rect -59 16 -55 17
rect -43 16 -39 32
<< ntransistor >>
rect -49 66 -45 68
rect -49 58 -45 60
rect -62 12 -60 16
rect -54 12 -52 16
<< ptransistor >>
rect -69 66 -65 68
rect -69 58 -65 60
rect -62 32 -60 36
rect -54 32 -52 36
<< ndcontact >>
rect -49 69 -45 73
rect -49 61 -45 65
rect -49 53 -45 57
rect -67 12 -63 16
rect -59 12 -55 16
rect -51 12 -47 16
<< pdcontact >>
rect -69 69 -65 73
rect -69 61 -65 65
rect -69 53 -65 57
rect -67 32 -63 36
rect -59 32 -55 36
rect -51 32 -47 36
<< m2contact >>
rect -69 77 -65 81
rect -49 77 -45 81
rect -76 61 -72 65
rect -64 61 -60 65
rect -54 61 -50 65
rect -69 45 -65 49
rect -49 45 -45 49
rect -59 37 -55 41
rect -75 32 -71 36
rect -43 32 -39 36
rect -59 27 -55 31
rect -59 17 -55 21
rect -75 12 -71 16
rect -43 12 -39 16
<< psubstratepcontact >>
rect -56 77 -52 81
rect -75 19 -71 23
rect -43 19 -39 23
<< nsubstratencontact >>
rect -62 45 -58 49
<< labels >>
rlabel polysilicon -62 6 -44 8 1 S0N
rlabel polysilicon -70 10 -68 40 1 S0
rlabel metal2 -75 16 -71 32 3 A
rlabel metal2 -43 16 -39 32 7 B
rlabel polysilicon -41 58 -39 76 7 S1N
rlabel metal2 -65 77 -49 81 5 C
rlabel polysilicon -73 50 -43 52 1 S1
rlabel m2contact -76 61 -72 65 3 OUT
<< end >>
