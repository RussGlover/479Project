magic
tech scmos
timestamp 1428433689
<< pwell >>
rect 11 -261 78 -244
rect 11 -329 36 -261
rect 66 -329 78 -261
rect 88 -310 142 -290
<< nwell >>
rect -5 -334 9 -309
rect 38 -334 64 -284
rect 80 -288 126 -276
rect 104 -324 150 -312
<< polysilicon >>
rect -4 -319 -2 -270
rect 89 -280 91 -263
rect 22 -295 28 -293
rect 32 -295 42 -293
rect 46 -295 52 -293
rect 22 -311 24 -295
rect 26 -299 28 -297
rect 32 -299 38 -297
rect 36 -301 38 -299
rect 50 -297 56 -295
rect 60 -297 70 -295
rect 74 -297 76 -295
rect 36 -303 42 -301
rect 46 -303 48 -301
rect 64 -301 70 -299
rect 74 -301 76 -299
rect 64 -303 66 -301
rect 36 -307 38 -303
rect 54 -305 56 -303
rect 60 -305 66 -303
rect 64 -307 66 -305
rect 89 -307 91 -284
rect 97 -290 99 -256
rect 115 -280 117 -263
rect 97 -292 112 -290
rect 97 -294 99 -292
rect 97 -300 99 -298
rect 110 -299 112 -292
rect 115 -297 117 -284
rect 123 -294 125 -256
rect 105 -302 107 -300
rect 110 -301 115 -299
rect 105 -307 107 -306
rect 64 -309 72 -307
rect 89 -309 107 -307
rect 70 -311 86 -309
rect 11 -313 24 -311
rect 84 -312 86 -311
rect 84 -314 95 -312
rect 64 -319 66 -316
rect 93 -316 95 -314
rect 113 -316 115 -301
rect 123 -312 125 -298
rect 131 -302 133 -263
rect 131 -308 133 -306
rect 123 -314 141 -312
rect 139 -316 141 -314
rect -4 -321 0 -319
rect 4 -321 14 -319
rect 18 -321 20 -319
rect 26 -321 28 -319
rect 32 -321 42 -319
rect 46 -321 50 -319
rect 54 -321 56 -319
rect 60 -321 70 -319
rect 74 -321 76 -319
rect 48 -327 50 -321
rect 113 -322 115 -320
rect 139 -322 141 -320
rect 127 -327 129 -324
rect 48 -328 84 -327
rect 98 -328 129 -327
rect 48 -329 129 -328
rect 82 -330 100 -329
<< ndiffusion >>
rect 28 -293 32 -292
rect 70 -295 74 -294
rect 28 -297 32 -295
rect 28 -300 32 -299
rect 70 -299 74 -297
rect 70 -302 74 -301
rect 96 -298 97 -294
rect 99 -298 100 -294
rect 122 -298 123 -294
rect 125 -298 126 -294
rect 104 -306 105 -302
rect 107 -306 108 -302
rect 14 -319 18 -318
rect 28 -319 32 -318
rect 70 -319 74 -318
rect 130 -306 131 -302
rect 133 -306 134 -302
rect 14 -322 18 -321
rect 28 -322 32 -321
rect 70 -322 74 -321
<< pdiffusion >>
rect 88 -284 89 -280
rect 91 -284 92 -280
rect 42 -293 46 -292
rect 56 -295 60 -294
rect 42 -296 46 -295
rect 42 -301 46 -300
rect 56 -298 60 -297
rect 56 -303 60 -302
rect 42 -304 46 -303
rect 56 -306 60 -305
rect 114 -284 115 -280
rect 117 -284 118 -280
rect 0 -319 4 -318
rect 42 -319 46 -318
rect 56 -319 60 -318
rect 112 -320 113 -316
rect 115 -320 116 -316
rect 138 -320 139 -316
rect 141 -320 142 -316
rect 0 -322 4 -321
rect 42 -322 46 -321
rect 56 -322 60 -321
<< metal1 >>
rect -14 -248 21 -244
rect 25 -248 50 -244
rect 56 -248 77 -244
rect 81 -248 150 -244
rect -14 -256 96 -252
rect 100 -256 122 -252
rect 126 -256 150 -252
rect -14 -263 88 -259
rect 92 -263 114 -259
rect 118 -263 130 -259
rect 134 -263 150 -259
rect -14 -270 -5 -266
rect -1 -270 150 -266
rect 70 -277 114 -273
rect 21 -288 25 -285
rect 35 -285 49 -281
rect 21 -292 28 -288
rect 4 -318 14 -314
rect 21 -322 25 -292
rect 35 -296 39 -285
rect 46 -290 53 -288
rect 70 -290 74 -277
rect 110 -280 114 -277
rect 46 -292 56 -290
rect 49 -294 56 -292
rect 63 -294 70 -290
rect 96 -284 104 -280
rect 84 -294 88 -284
rect 100 -294 104 -284
rect 35 -300 42 -296
rect 32 -304 39 -300
rect 49 -304 53 -294
rect 63 -298 67 -294
rect 60 -302 67 -298
rect 84 -298 92 -294
rect 122 -284 130 -280
rect 110 -294 114 -284
rect 126 -294 130 -284
rect 110 -298 118 -294
rect 32 -311 35 -307
rect 46 -306 53 -304
rect 46 -308 56 -306
rect 35 -314 39 -311
rect 49 -310 56 -308
rect 49 -314 53 -310
rect 63 -312 67 -302
rect 74 -306 77 -302
rect 32 -318 42 -314
rect 49 -318 56 -314
rect 74 -318 76 -314
rect 49 -322 53 -318
rect 84 -322 88 -298
rect 100 -302 104 -298
rect 126 -302 130 -298
rect 112 -306 120 -302
rect 100 -316 104 -306
rect 116 -316 120 -306
rect 97 -320 108 -316
rect 18 -326 28 -322
rect 46 -326 53 -322
rect 60 -326 70 -322
rect 74 -326 88 -322
rect 116 -323 120 -320
rect 0 -330 4 -326
rect 49 -330 53 -326
rect 96 -327 120 -323
rect 138 -306 146 -302
rect 126 -316 130 -306
rect 142 -316 146 -306
rect 126 -320 134 -316
rect 142 -323 146 -320
rect -14 -334 -1 -330
rect 5 -334 48 -330
rect 54 -334 150 -330
<< metal2 >>
rect 21 -281 25 -248
rect 24 -324 28 -307
rect 17 -328 28 -324
rect 17 -334 21 -328
rect 40 -334 44 -244
rect 49 -323 53 -285
rect 77 -302 81 -248
rect 76 -306 77 -302
rect 76 -311 81 -306
rect 76 -314 80 -311
rect 84 -319 104 -315
rect 84 -323 88 -319
rect 100 -323 104 -319
rect 49 -327 88 -323
rect 100 -327 142 -323
rect 92 -334 96 -327
<< ntransistor >>
rect 28 -295 32 -293
rect 28 -299 32 -297
rect 70 -297 74 -295
rect 70 -301 74 -299
rect 97 -298 99 -294
rect 123 -298 125 -294
rect 105 -306 107 -302
rect 131 -306 133 -302
rect 14 -321 18 -319
rect 28 -321 32 -319
rect 70 -321 74 -319
<< ptransistor >>
rect 89 -284 91 -280
rect 42 -295 46 -293
rect 56 -297 60 -295
rect 42 -303 46 -301
rect 56 -305 60 -303
rect 115 -284 117 -280
rect 0 -321 4 -319
rect 42 -321 46 -319
rect 56 -321 60 -319
rect 113 -320 115 -316
rect 139 -320 141 -316
<< polycontact >>
rect 96 -256 100 -252
rect 122 -256 126 -252
rect 88 -263 92 -259
rect -5 -270 -1 -266
rect 7 -314 11 -310
rect 35 -311 39 -307
rect 114 -263 118 -259
rect 130 -263 134 -259
rect 63 -316 67 -312
rect 93 -320 97 -316
rect 126 -324 130 -320
<< ndcontact >>
rect 28 -292 32 -288
rect 70 -294 74 -290
rect 28 -304 32 -300
rect 70 -306 74 -302
rect 92 -298 96 -294
rect 100 -298 104 -294
rect 118 -298 122 -294
rect 126 -298 130 -294
rect 100 -306 104 -302
rect 108 -306 112 -302
rect 14 -318 18 -314
rect 28 -318 32 -314
rect 70 -318 74 -314
rect 126 -306 130 -302
rect 134 -306 138 -302
rect 14 -326 18 -322
rect 28 -326 32 -322
rect 70 -326 74 -322
<< pdcontact >>
rect 84 -284 88 -280
rect 92 -284 96 -280
rect 42 -292 46 -288
rect 56 -294 60 -290
rect 42 -300 46 -296
rect 56 -302 60 -298
rect 42 -308 46 -304
rect 56 -310 60 -306
rect 110 -284 114 -280
rect 118 -284 122 -280
rect 0 -318 4 -314
rect 42 -318 46 -314
rect 56 -318 60 -314
rect 108 -320 112 -316
rect 116 -320 120 -316
rect 134 -320 138 -316
rect 142 -320 146 -316
rect 0 -326 4 -322
rect 42 -326 46 -322
rect 56 -326 60 -322
<< m2contact >>
rect 21 -248 25 -244
rect 77 -248 81 -244
rect 21 -285 25 -281
rect 49 -285 53 -281
rect 28 -311 32 -307
rect 77 -306 81 -302
rect 76 -318 80 -314
rect 92 -327 96 -323
rect 142 -327 146 -323
<< psubstratepcontact >>
rect 50 -248 56 -244
<< nsubstratencontact >>
rect -1 -334 5 -330
rect 48 -334 54 -330
<< labels >>
rlabel metal1 148 -332 148 -332 8 Vdd
rlabel metal2 19 -332 19 -332 1 Q
rlabel metal2 42 -332 42 -332 1 dividendin
rlabel metal2 94 -332 94 -332 1 D
rlabel metal1 148 -268 148 -268 7 rst
rlabel metal1 148 -261 148 -261 7 CB
rlabel metal1 148 -254 148 -254 7 C
rlabel metal1 148 -246 148 -246 7 GND
<< end >>
