magic
tech scmos
timestamp 1428666073
<< nwell >>
rect -65 25 -47 36
rect -114 -35 88 9
<< polysilicon >>
rect -47 57 -45 59
rect -26 57 31 59
rect -103 49 -101 51
rect -75 49 -73 51
rect -47 49 -45 53
rect -36 49 -34 51
rect -26 49 -24 57
rect -22 53 21 55
rect -22 49 -20 53
rect -18 49 -16 51
rect -1 49 1 51
rect 8 49 10 51
rect 19 49 21 53
rect 29 49 31 57
rect 39 57 79 59
rect 39 49 41 57
rect 43 53 67 55
rect 43 49 45 53
rect 54 49 56 51
rect 65 49 67 53
rect 77 49 79 57
rect -103 6 -101 43
rect -103 -12 -101 2
rect -75 -6 -73 43
rect -47 38 -45 43
rect -57 36 -45 38
rect -57 33 -55 36
rect -57 26 -55 29
rect -36 24 -34 43
rect -75 -12 -73 -10
rect -36 -12 -34 20
rect -26 -12 -24 43
rect -22 -12 -20 43
rect -18 8 -16 43
rect -1 15 1 43
rect 8 9 10 43
rect 19 37 21 43
rect 29 41 31 43
rect 39 41 41 43
rect 29 39 41 41
rect 43 37 45 43
rect 19 35 45 37
rect 40 34 44 35
rect 54 10 56 43
rect -18 6 8 8
rect -18 -12 -16 6
rect -1 -12 1 -2
rect 8 -12 10 5
rect 19 -6 45 -4
rect 19 -12 21 -6
rect 29 -10 41 -8
rect 29 -12 31 -10
rect 39 -12 41 -10
rect 43 -12 45 -6
rect 54 -12 56 6
rect 65 -12 67 43
rect 77 41 79 43
rect 77 -3 81 -1
rect 77 -12 79 -3
rect -103 -20 -101 -18
rect -75 -20 -73 -18
rect -36 -20 -34 -18
rect -26 -26 -24 -18
rect -22 -22 -20 -18
rect -18 -20 -16 -18
rect -1 -20 1 -18
rect 8 -20 10 -18
rect 19 -22 21 -18
rect -22 -24 21 -22
rect 29 -26 31 -18
rect -26 -28 31 -26
rect 39 -26 41 -18
rect 43 -22 45 -18
rect 54 -20 56 -18
rect 65 -22 67 -18
rect 43 -24 67 -22
rect 77 -26 79 -18
rect 39 -28 79 -26
<< ndiffusion >>
rect -114 48 -103 49
rect -114 43 -111 48
rect -107 43 -103 48
rect -101 48 -93 49
rect -101 44 -99 48
rect -95 44 -93 48
rect -101 43 -93 44
rect -87 48 -75 49
rect -87 44 -83 48
rect -79 44 -75 48
rect -87 43 -75 44
rect -73 48 -65 49
rect -73 44 -71 48
rect -67 44 -65 48
rect -73 43 -65 44
rect -62 48 -47 49
rect -62 44 -53 48
rect -49 44 -47 48
rect -62 43 -47 44
rect -45 48 -36 49
rect -45 44 -42 48
rect -38 44 -36 48
rect -45 43 -36 44
rect -34 48 -26 49
rect -34 44 -32 48
rect -28 44 -26 48
rect -34 43 -26 44
rect -24 43 -22 49
rect -20 43 -18 49
rect -16 48 -1 49
rect -16 44 -11 48
rect -7 44 -1 48
rect -16 43 -1 44
rect 1 48 8 49
rect 1 44 2 48
rect 6 44 8 48
rect 1 43 8 44
rect 10 48 19 49
rect 10 44 12 48
rect 16 44 19 48
rect 10 43 19 44
rect 21 48 29 49
rect 21 44 23 48
rect 27 44 29 48
rect 21 43 29 44
rect 31 48 39 49
rect 31 44 33 48
rect 37 44 39 48
rect 31 43 39 44
rect 41 43 43 49
rect 45 48 54 49
rect 45 44 47 48
rect 51 44 54 48
rect 45 43 54 44
rect 56 48 65 49
rect 56 44 58 48
rect 62 44 65 48
rect 56 43 65 44
rect 67 48 77 49
rect 67 44 69 48
rect 73 44 77 48
rect 67 43 77 44
rect 79 48 88 49
rect 79 44 82 48
rect 86 44 88 48
rect 79 43 88 44
<< pdiffusion >>
rect -59 29 -57 33
rect -55 29 -53 33
rect -114 -13 -103 -12
rect -114 -17 -111 -13
rect -107 -17 -103 -13
rect -114 -18 -103 -17
rect -101 -13 -93 -12
rect -101 -17 -99 -13
rect -95 -17 -93 -13
rect -101 -18 -93 -17
rect -87 -13 -75 -12
rect -87 -17 -83 -13
rect -79 -17 -75 -13
rect -87 -18 -75 -17
rect -73 -13 -65 -12
rect -73 -17 -71 -13
rect -67 -17 -65 -13
rect -73 -18 -65 -17
rect -45 -13 -36 -12
rect -45 -17 -42 -13
rect -38 -17 -36 -13
rect -45 -18 -36 -17
rect -34 -13 -26 -12
rect -34 -17 -32 -13
rect -28 -17 -26 -13
rect -34 -18 -26 -17
rect -24 -18 -22 -12
rect -20 -18 -18 -12
rect -16 -13 -1 -12
rect -16 -17 -11 -13
rect -7 -17 -1 -13
rect -16 -18 -1 -17
rect 1 -13 8 -12
rect 1 -17 2 -13
rect 6 -17 8 -13
rect 1 -18 8 -17
rect 10 -13 19 -12
rect 10 -17 12 -13
rect 16 -17 19 -13
rect 10 -18 19 -17
rect 21 -13 29 -12
rect 21 -17 23 -13
rect 27 -17 29 -13
rect 21 -18 29 -17
rect 31 -13 39 -12
rect 31 -17 33 -13
rect 37 -17 39 -13
rect 31 -18 39 -17
rect 41 -18 43 -12
rect 45 -13 54 -12
rect 45 -17 47 -13
rect 51 -17 54 -13
rect 45 -18 54 -17
rect 56 -13 65 -12
rect 56 -17 58 -13
rect 62 -17 65 -13
rect 56 -18 65 -17
rect 67 -13 77 -12
rect 67 -18 70 -13
rect 74 -18 77 -13
rect 79 -13 88 -12
rect 79 -17 82 -13
rect 86 -17 88 -13
rect 79 -18 88 -17
<< metal1 >>
rect -132 75 -128 79
rect 6 75 19 79
rect 12 65 16 75
rect -114 61 97 65
rect -99 48 -95 61
rect -71 48 -67 61
rect -43 53 -39 57
rect -32 48 -28 61
rect 12 48 16 61
rect 33 48 37 61
rect 69 48 73 61
rect -111 40 -107 44
rect -83 37 -79 44
rect -53 33 -49 44
rect -42 40 -38 44
rect -11 40 -7 44
rect 2 41 6 44
rect 23 41 27 44
rect 2 37 27 41
rect 47 39 51 44
rect 58 40 62 44
rect 82 40 86 44
rect 58 36 86 40
rect -4 33 40 34
rect -49 30 40 33
rect -49 29 -2 30
rect -63 24 -59 29
rect -116 20 -38 24
rect -34 20 96 24
rect -46 10 -32 14
rect 3 12 39 16
rect 3 11 5 12
rect -116 6 -111 10
rect -1 6 3 11
rect 47 9 52 10
rect -100 2 3 6
rect 12 6 52 9
rect 56 6 96 10
rect 12 5 48 6
rect 3 -2 51 2
rect 62 -1 77 3
rect -111 -13 -107 -9
rect -83 -13 -79 -6
rect -71 -10 -50 -6
rect -42 -13 -38 -9
rect -28 -10 -11 -6
rect -11 -13 -7 -10
rect 2 -10 27 -6
rect 2 -13 6 -10
rect 23 -13 27 -10
rect 47 -13 51 -2
rect 58 -9 86 -5
rect 58 -13 62 -9
rect 82 -13 86 -9
rect -99 -31 -95 -17
rect -71 -31 -67 -17
rect -32 -31 -28 -17
rect 12 -31 16 -17
rect 33 -31 37 -17
rect 70 -31 74 -17
rect -114 -35 88 -31
<< metal2 >>
rect -33 57 -29 71
rect -48 53 -43 57
rect -35 53 -29 57
rect -111 10 -107 36
rect -111 -5 -107 6
rect -83 -2 -79 33
rect -83 -44 -79 -6
rect -50 -6 -46 10
rect -42 -5 -38 36
rect -32 -6 -28 10
rect -22 -43 -18 71
rect -11 -6 -7 36
rect -1 -2 3 2
rect 30 -39 34 69
rect 47 16 51 35
rect 43 12 51 16
rect 58 3 62 71
<< ntransistor >>
rect -103 43 -101 49
rect -75 43 -73 49
rect -47 43 -45 49
rect -36 43 -34 49
rect -26 43 -24 49
rect -22 43 -20 49
rect -18 43 -16 49
rect -1 43 1 49
rect 8 43 10 49
rect 19 43 21 49
rect 29 43 31 49
rect 39 43 41 49
rect 43 43 45 49
rect 54 43 56 49
rect 65 43 67 49
rect 77 43 79 49
<< ptransistor >>
rect -57 29 -55 33
rect -103 -18 -101 -12
rect -75 -18 -73 -12
rect -36 -18 -34 -12
rect -26 -18 -24 -12
rect -22 -18 -20 -12
rect -18 -18 -16 -12
rect -1 -18 1 -12
rect 8 -18 10 -12
rect 19 -18 21 -12
rect 29 -18 31 -12
rect 39 -18 41 -12
rect 43 -18 45 -12
rect 54 -18 56 -12
rect 65 -18 67 -12
rect 77 -18 79 -12
<< polycontact >>
rect -47 53 -43 57
rect -104 2 -100 6
rect -38 20 -34 24
rect -75 -10 -71 -6
rect -1 11 3 15
rect 40 30 44 34
rect 8 5 12 9
rect 52 6 56 10
rect -1 -2 3 2
rect 77 -1 81 3
<< ndcontact >>
rect -111 44 -107 48
rect -99 44 -95 48
rect -83 44 -79 48
rect -71 44 -67 48
rect -53 44 -49 48
rect -42 44 -38 48
rect -32 44 -28 48
rect -11 44 -7 48
rect 2 44 6 48
rect 12 44 16 48
rect 23 44 27 48
rect 33 44 37 48
rect 47 44 51 48
rect 58 44 62 48
rect 69 44 73 48
rect 82 44 86 48
<< pdcontact >>
rect -63 29 -59 33
rect -53 29 -49 33
rect -111 -17 -107 -13
rect -99 -17 -95 -13
rect -83 -17 -79 -13
rect -71 -17 -67 -13
rect -42 -17 -38 -13
rect -32 -17 -28 -13
rect -11 -17 -7 -13
rect 2 -17 6 -13
rect 12 -17 16 -13
rect 23 -17 27 -13
rect 33 -17 37 -13
rect 47 -17 51 -13
rect 58 -17 62 -13
rect 70 -17 74 -13
rect 82 -17 86 -13
<< m2contact >>
rect -39 53 -35 57
rect -111 36 -107 40
rect -83 33 -79 37
rect -42 36 -38 40
rect -11 36 -7 40
rect 47 35 51 39
rect -50 10 -46 14
rect -32 10 -28 14
rect 39 12 43 16
rect -111 6 -107 10
rect 58 -1 62 3
rect -111 -9 -107 -5
rect -83 -6 -79 -2
rect -50 -10 -46 -6
rect -42 -9 -38 -5
rect -32 -10 -28 -6
rect -11 -10 -7 -6
<< labels >>
rlabel metal2 -33 71 -29 71 5 B
rlabel metal2 30 69 34 69 5 fromShift
rlabel metal2 -83 -44 -79 -44 1 Z
rlabel metal1 -116 6 -116 10 3 x
rlabel metal1 96 20 96 24 7 Add
rlabel metal2 58 71 62 71 1 A
rlabel metal1 -114 61 -114 65 1 Gnd
rlabel metal1 -114 -35 -114 -31 1 Vdd
rlabel metal1 96 6 96 10 7 C
rlabel metal1 -31 29 -31 33 1 xor
<< end >>
