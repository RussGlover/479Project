magic
tech scmos
timestamp 1428802636
<< metal1 >>
rect 65 4 74 8
rect 65 -18 74 -14
rect 65 -25 74 -21
rect 65 -32 74 -28
rect 65 -158 74 -154
use reg11  reg11_0
timestamp 1428636301
transform 1 0 96 0 1 18
box -113 -176 -31 -10
use reg11  reg11_1
timestamp 1428636301
transform 1 0 187 0 1 18
box -113 -176 -31 -10
<< end >>
