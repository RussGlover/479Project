magic
tech scmos
timestamp 1428734395
<< metal1 >>
rect 166 159 175 163
rect 166 151 175 155
rect 166 144 175 148
rect 166 137 175 141
rect 166 130 175 134
rect 166 123 175 127
rect 166 -3 175 1
rect 166 -17 175 -13
rect 166 -71 175 -67
rect 166 -85 175 -81
rect 156 -126 175 -122
rect 165 -134 175 -130
rect 165 -143 175 -139
rect 71 -151 127 -147
rect 127 -161 131 -157
rect 165 -161 175 -157
rect 165 -180 175 -176
rect 159 -192 175 -188
rect 159 -199 175 -195
rect 159 -218 175 -214
rect 159 -225 175 -221
rect 159 -232 175 -228
<< metal2 >>
rect -3 163 1 166
rect 47 159 51 166
rect 36 -7 40 -2
rect 47 -8 51 -3
rect 108 -5 112 -3
rect 99 -9 112 -5
rect 127 -7 131 -3
rect 127 -147 131 -55
rect 127 -212 131 -151
<< m2contact >>
rect 127 -151 131 -147
use reg1  reg1_0
timestamp 1428711541
transform 1 0 106 0 1 173
box -144 -176 -18 -10
use rr1  rr1_0
timestamp 1428723998
transform 1 0 197 0 1 173
box -113 -176 -31 -10
use mux1  mux1_0
timestamp 1428729551
transform 1 0 102 0 1 -161
box -140 -27 64 31
use dp1v2  shift1_0
timestamp 1428712110
transform 1 0 11 0 1 -12
box -49 -220 155 13
<< labels >>
rlabel metal2 47 166 51 166 5 dividendin
rlabel metal2 -3 166 1 166 5 divisorin
rlabel metal1 169 159 169 163 6 Vdd
rlabel metal1 169 151 169 155 7 clockload
rlabel metal1 169 144 169 148 7 notclockload
rlabel metal1 169 137 169 141 7 clk
rlabel metal1 169 130 169 134 7 notclk
rlabel metal1 169 123 169 127 7 reset
rlabel metal2 127 -212 131 -212 1 remainder
rlabel metal1 169 -17 169 -13 7 Gnd
rlabel metal1 162 -192 162 -188 1 Gnd
rlabel metal1 162 -199 162 -195 1 inbit
rlabel metal1 162 -218 162 -214 1 notshift
rlabel metal1 162 -225 162 -221 1 shift
rlabel metal1 162 -232 162 -228 1 Vdd
rlabel metal1 170 -126 170 -122 7 Vdd
rlabel metal1 175 -71 175 -67 7 Add
rlabel metal1 175 -85 175 -81 7 C
rlabel metal1 171 -134 171 -130 7 S1n
rlabel metal1 171 -143 171 -139 7 S0n
rlabel metal1 171 -161 171 -157 7 S0
rlabel metal1 171 -180 171 -176 7 S1
<< end >>
