magic
tech scmos
timestamp 1428985832
<< metal1 >>
rect 166 159 175 163
rect 166 151 175 155
rect 166 144 175 148
rect 166 137 175 141
rect 166 130 175 134
rect 166 123 175 127
rect 166 -3 175 1
rect 166 -17 175 -13
rect 166 -71 175 -67
rect 166 -85 175 -81
rect 156 -126 175 -122
rect 165 -134 175 -130
rect 165 -143 175 -139
rect 127 -161 131 -157
rect 165 -161 175 -157
rect 165 -180 175 -176
rect 159 -192 175 -188
rect 159 -199 175 -195
rect 159 -218 175 -214
rect 159 -225 175 -221
rect 159 -232 175 -228
<< metal2 >>
rect -3 163 1 166
rect 47 159 51 166
rect 36 -7 40 -2
rect 47 -8 51 -3
rect 108 -5 112 -3
rect 99 -9 112 -5
rect 127 -7 131 -3
rect 127 -147 131 -55
rect 127 -212 131 -151
<< m2contact >>
rect 127 -151 131 -147
use reg1  reg1_0
timestamp 1428981317
transform 1 0 106 0 1 173
box -144 -176 -18 -10
use rr1  rr1_0
timestamp 1428973229
transform 1 0 197 0 1 173
box -113 -176 -31 -10
use mux1  mux1_0
timestamp 1428963193
transform 1 0 102 0 1 -161
box -140 -31 64 31
use dp1v2  shift1_0
timestamp 1428973275
transform 1 0 11 0 1 -12
box -49 -220 155 13
<< end >>
