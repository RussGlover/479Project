magic
tech scmos
timestamp 1428734601
<< metal1 >>
rect 145 87 182 91
rect 145 79 182 83
rect 145 72 182 76
rect 145 65 182 69
rect 145 58 182 62
rect 145 51 182 55
rect 17 -190 106 -186
rect 87 -223 143 -219
rect -22 -264 -18 -260
rect 145 -264 182 -260
rect -22 -271 -18 -267
rect 145 -271 182 -267
rect -22 -290 -18 -286
rect 145 -290 182 -286
rect -22 -297 -18 -293
rect 145 -297 182 -293
rect -22 -304 -18 -300
rect 145 -304 182 -300
<< metal2 >>
rect 13 -207 17 -190
rect 46 -202 50 95
rect 87 -195 91 -75
rect 106 -186 110 -70
rect 110 -190 147 -186
rect 87 -199 107 -195
rect 103 -256 107 -199
rect 143 -200 147 -190
rect 88 -260 107 -256
<< m2contact >>
rect 13 -190 17 -186
rect 106 -190 110 -186
rect 143 -223 147 -219
use rr1  rr1_0
timestamp 1428723998
transform 1 0 176 0 1 101
box -113 -176 -31 -10
use mux1  mux1_0
timestamp 1428729551
transform 1 0 118 0 1 -233
box -140 -27 64 31
use shift1  shift1_0
timestamp 1428723798
transform 1 0 0 0 1 -108
box -18 -196 146 -152
<< end >>
