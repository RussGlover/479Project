magic
tech scmos
timestamp 1428369478
<< pwell >>
rect -113 -102 -85 -76
rect -113 -158 -85 -132
rect -47 -176 -31 -54
<< nwell >>
rect -82 -62 -49 -10
rect -113 -74 -49 -62
rect -74 -104 -49 -74
rect -113 -130 -49 -104
rect -74 -160 -49 -130
rect -113 -176 -49 -160
<< polysilicon >>
rect -102 -63 -100 -36
rect -104 -65 -100 -63
rect -104 -66 -102 -65
rect -104 -94 -102 -70
rect -96 -80 -94 -43
rect -89 -63 -87 -50
rect -46 -56 -33 -54
rect -89 -65 -57 -63
rect -53 -65 -43 -63
rect -39 -65 -37 -63
rect -35 -79 -33 -56
rect -104 -122 -102 -98
rect -96 -108 -94 -84
rect -86 -87 -84 -79
rect -59 -81 -57 -79
rect -53 -81 -43 -79
rect -39 -81 -33 -79
rect -48 -85 -43 -83
rect -39 -85 -37 -83
rect -48 -87 -46 -85
rect -86 -89 -57 -87
rect -53 -89 -46 -87
rect -65 -111 -57 -109
rect -53 -111 -43 -109
rect -39 -111 -37 -109
rect -104 -150 -102 -126
rect -96 -136 -94 -112
rect -65 -136 -63 -111
rect -35 -131 -33 -81
rect -59 -133 -57 -131
rect -53 -133 -42 -131
rect -38 -133 -33 -131
rect -74 -138 -63 -136
rect -49 -137 -42 -135
rect -38 -137 -36 -135
rect -49 -139 -47 -137
rect -104 -156 -102 -154
rect -96 -164 -94 -140
rect -61 -141 -57 -139
rect -53 -141 -47 -139
rect -87 -146 -73 -144
rect -49 -146 -47 -141
rect -75 -152 -73 -146
rect -75 -154 -61 -152
rect -63 -155 -61 -154
rect -63 -157 -57 -155
rect -53 -157 -43 -155
rect -39 -157 -37 -155
rect -96 -170 -94 -168
<< ndiffusion >>
rect -43 -63 -39 -62
rect -43 -66 -39 -65
rect -43 -79 -39 -78
rect -97 -84 -96 -80
rect -94 -84 -93 -80
rect -105 -98 -104 -94
rect -102 -98 -101 -94
rect -43 -83 -39 -81
rect -43 -86 -39 -85
rect -43 -109 -39 -108
rect -97 -140 -96 -136
rect -94 -140 -93 -136
rect -43 -112 -39 -111
rect -42 -131 -38 -130
rect -42 -135 -38 -133
rect -105 -154 -104 -150
rect -102 -154 -101 -150
rect -42 -138 -38 -137
rect -43 -155 -39 -154
rect -43 -158 -39 -157
<< pdiffusion >>
rect -105 -70 -104 -66
rect -102 -70 -101 -66
rect -57 -63 -53 -62
rect -57 -66 -53 -65
rect -57 -79 -53 -78
rect -57 -82 -53 -81
rect -57 -87 -53 -86
rect -57 -90 -53 -89
rect -97 -112 -96 -108
rect -94 -112 -93 -108
rect -57 -109 -53 -108
rect -105 -126 -104 -122
rect -102 -126 -101 -122
rect -57 -112 -53 -111
rect -57 -131 -53 -130
rect -57 -134 -53 -133
rect -57 -139 -53 -138
rect -57 -142 -53 -141
rect -57 -155 -53 -154
rect -57 -158 -53 -157
rect -97 -168 -96 -164
rect -94 -168 -93 -164
<< metal1 >>
rect -113 -14 -79 -10
rect -73 -14 -70 -10
rect -66 -14 -31 -10
rect -113 -22 -31 -18
rect -113 -29 -31 -25
rect -113 -36 -103 -32
rect -99 -36 -31 -32
rect -113 -43 -97 -39
rect -93 -43 -31 -39
rect -113 -50 -90 -46
rect -86 -50 -31 -46
rect -50 -58 -46 -57
rect -53 -62 -43 -58
rect -109 -66 -105 -65
rect -97 -70 -89 -66
rect -66 -70 -57 -66
rect -39 -70 -31 -66
rect -109 -80 -105 -70
rect -93 -75 -89 -70
rect -93 -79 -87 -75
rect -66 -78 -57 -74
rect -50 -78 -43 -74
rect -93 -80 -89 -79
rect -109 -84 -101 -80
rect -50 -82 -46 -78
rect -93 -87 -89 -84
rect -53 -86 -46 -82
rect -35 -86 -31 -70
rect -109 -91 -89 -87
rect -109 -94 -105 -91
rect -66 -94 -57 -90
rect -97 -98 -89 -94
rect -50 -97 -46 -86
rect -39 -90 -31 -86
rect -109 -108 -105 -98
rect -93 -104 -89 -98
rect -74 -101 -46 -97
rect -93 -108 -57 -104
rect -53 -108 -43 -104
rect -109 -112 -101 -108
rect -35 -112 -31 -90
rect -109 -119 -82 -115
rect -66 -116 -57 -112
rect -39 -116 -31 -112
rect -109 -122 -105 -119
rect -97 -126 -89 -122
rect -86 -123 -45 -119
rect -49 -126 -45 -123
rect -109 -136 -105 -126
rect -93 -136 -89 -126
rect -66 -130 -57 -126
rect -49 -130 -42 -126
rect -109 -140 -101 -136
rect -93 -143 -89 -140
rect -49 -134 -45 -130
rect -78 -135 -74 -134
rect -53 -138 -45 -134
rect -35 -138 -31 -116
rect -109 -147 -91 -143
rect -109 -150 -105 -147
rect -78 -150 -74 -139
rect -38 -142 -31 -138
rect -66 -146 -57 -142
rect -97 -154 -74 -150
rect -53 -154 -43 -150
rect -109 -164 -105 -154
rect -93 -164 -89 -154
rect -66 -159 -57 -158
rect -70 -162 -57 -159
rect -109 -168 -101 -164
rect -50 -165 -46 -154
rect -35 -158 -31 -142
rect -39 -162 -31 -158
rect -66 -169 -46 -165
rect -113 -176 -41 -172
rect -35 -176 -31 -162
<< metal2 >>
rect -109 -61 -85 -57
rect -89 -176 -85 -61
rect -70 -66 -66 -14
rect -70 -74 -66 -70
rect -70 -90 -66 -78
rect -78 -130 -74 -101
rect -70 -112 -66 -94
rect -70 -126 -66 -116
rect -70 -142 -66 -130
rect -70 -155 -66 -146
rect -70 -176 -66 -169
<< ntransistor >>
rect -43 -65 -39 -63
rect -96 -84 -94 -80
rect -104 -98 -102 -94
rect -43 -81 -39 -79
rect -43 -85 -39 -83
rect -43 -111 -39 -109
rect -96 -140 -94 -136
rect -42 -133 -38 -131
rect -42 -137 -38 -135
rect -104 -154 -102 -150
rect -43 -157 -39 -155
<< ptransistor >>
rect -104 -70 -102 -66
rect -57 -65 -53 -63
rect -57 -81 -53 -79
rect -57 -89 -53 -87
rect -96 -112 -94 -108
rect -57 -111 -53 -109
rect -104 -126 -102 -122
rect -57 -133 -53 -131
rect -57 -141 -53 -139
rect -57 -157 -53 -155
rect -96 -168 -94 -164
<< polycontact >>
rect -103 -36 -99 -32
rect -97 -43 -93 -39
rect -90 -50 -86 -46
rect -50 -57 -46 -53
rect -87 -79 -83 -75
rect -78 -139 -74 -135
rect -91 -147 -87 -143
rect -50 -150 -46 -146
<< ndcontact >>
rect -43 -62 -39 -58
rect -43 -70 -39 -66
rect -43 -78 -39 -74
rect -101 -84 -97 -80
rect -93 -84 -89 -80
rect -109 -98 -105 -94
rect -101 -98 -97 -94
rect -43 -90 -39 -86
rect -43 -108 -39 -104
rect -101 -140 -97 -136
rect -93 -140 -89 -136
rect -43 -116 -39 -112
rect -42 -130 -38 -126
rect -109 -154 -105 -150
rect -101 -154 -97 -150
rect -42 -142 -38 -138
rect -43 -154 -39 -150
rect -43 -162 -39 -158
<< pdcontact >>
rect -109 -70 -105 -66
rect -101 -70 -97 -66
rect -57 -62 -53 -58
rect -57 -70 -53 -66
rect -57 -78 -53 -74
rect -57 -86 -53 -82
rect -57 -94 -53 -90
rect -57 -108 -53 -104
rect -101 -112 -97 -108
rect -93 -112 -89 -108
rect -109 -126 -105 -122
rect -101 -126 -97 -122
rect -57 -116 -53 -112
rect -57 -130 -53 -126
rect -57 -138 -53 -134
rect -57 -146 -53 -142
rect -57 -154 -53 -150
rect -57 -162 -53 -158
rect -101 -168 -97 -164
rect -93 -168 -89 -164
<< m2contact >>
rect -70 -14 -66 -10
rect -109 -65 -105 -61
rect -70 -70 -66 -66
rect -70 -78 -66 -74
rect -70 -94 -66 -90
rect -78 -101 -74 -97
rect -70 -116 -66 -112
rect -70 -130 -66 -126
rect -78 -134 -74 -130
rect -70 -146 -66 -142
rect -70 -159 -66 -155
rect -70 -169 -66 -165
<< psubstratepcontact >>
rect -41 -176 -35 -172
<< nsubstratencontact >>
rect -79 -14 -73 -10
<< labels >>
rlabel metal2 -68 -174 -68 -174 1 Q
rlabel metal1 -33 -174 -33 -174 1 GND
rlabel metal1 -33 -12 -33 -12 7 Vdd
rlabel metal1 -33 -48 -33 -48 7 rst
rlabel metal1 -33 -41 -33 -41 7 CB
rlabel metal1 -33 -34 -33 -34 7 C
rlabel metal2 -87 -174 -87 -174 1 D
rlabel metal1 -33 -20 -33 -20 7 Cl
rlabel metal1 -33 -27 -33 -27 7 ClB
<< end >>
