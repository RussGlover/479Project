magic
tech scmos
timestamp 1428565332
<< metal2 >>
rect 36 -7 40 -2
rect 47 -8 51 -3
rect 108 -5 112 -3
rect 99 -9 112 -5
rect 127 -7 131 -3
rect 103 -106 110 -102
rect 106 -160 110 -106
rect 99 -164 110 -160
use reg1  reg1_0
timestamp 1428364277
transform 1 0 106 0 1 173
box -113 -176 -31 -23
use rr1  rr1_0
timestamp 1428369478
transform 1 0 197 0 1 173
box -113 -176 -31 -10
use adder7  adder7_0
timestamp 1428559628
transform 1 0 69 0 1 -78
box -78 -33 97 79
use mux1  mux1_0
timestamp 1428565219
transform 1 0 102 0 1 -161
box -82 -3 29 93
use shift1  shift1_0
timestamp 1428367300
transform 1 0 11 0 1 -12
box -18 -196 146 -152
<< end >>
