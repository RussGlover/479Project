magic
tech scmos
timestamp 1428973275
<< pwell >>
rect -10 -202 84 -176
rect -10 -214 17 -202
<< nwell >>
rect 28 -220 98 -206
<< polysilicon >>
rect 0 -185 78 -183
rect 0 -195 2 -185
rect -20 -197 -6 -195
rect -2 -197 2 -195
rect 4 -189 72 -187
rect 4 -203 6 -189
rect 38 -195 40 -193
rect 58 -195 60 -193
rect 14 -201 21 -199
rect 19 -202 21 -201
rect 38 -202 40 -199
rect -11 -205 -6 -203
rect -2 -205 6 -203
rect 19 -204 40 -202
rect 38 -209 40 -204
rect 58 -203 60 -199
rect 47 -205 60 -203
rect 58 -209 60 -205
rect 70 -209 72 -189
rect 76 -202 78 -185
rect 38 -215 40 -213
rect 58 -215 60 -213
<< ndiffusion >>
rect -6 -195 -2 -194
rect -6 -198 -2 -197
rect -6 -203 -2 -202
rect 37 -199 38 -195
rect 40 -199 41 -195
rect 57 -199 58 -195
rect 60 -199 61 -195
rect -6 -206 -2 -205
<< pdiffusion >>
rect 37 -213 38 -209
rect 40 -213 41 -209
rect 57 -213 58 -209
rect 60 -213 61 -209
<< metal1 >>
rect 94 -139 118 -135
rect -49 -180 28 -176
rect 32 -180 34 -176
rect 46 -180 48 -176
rect 52 -180 150 -176
rect -49 -187 -6 -183
rect -6 -190 -2 -187
rect 18 -187 149 -183
rect 18 -192 22 -187
rect 65 -194 101 -190
rect 61 -195 65 -194
rect -24 -202 -20 -198
rect -2 -202 10 -198
rect 32 -199 33 -195
rect 52 -199 53 -195
rect 41 -202 45 -199
rect -49 -206 -20 -202
rect 41 -206 43 -202
rect -15 -209 -11 -206
rect -49 -213 -11 -209
rect -2 -210 18 -206
rect 41 -209 45 -206
rect 61 -209 65 -199
rect 79 -206 148 -202
rect 73 -213 148 -209
rect 33 -216 37 -213
rect 53 -216 57 -213
rect -49 -220 79 -216
rect 91 -220 148 -216
<< metal2 >>
rect 92 -118 105 -114
rect 71 -176 90 -172
rect 1 -183 5 -176
rect -2 -187 5 -183
rect 1 -214 5 -187
rect 18 -206 22 -196
rect 28 -195 32 -180
rect 48 -195 52 -180
rect 86 -214 90 -176
rect 101 -190 105 -118
rect 1 -218 90 -214
<< ntransistor >>
rect -6 -197 -2 -195
rect 38 -199 40 -195
rect 58 -199 60 -195
rect -6 -205 -2 -203
<< ptransistor >>
rect 38 -213 40 -209
rect 58 -213 60 -209
<< polycontact >>
rect -24 -198 -20 -194
rect -15 -206 -11 -202
rect 10 -202 14 -198
rect 43 -206 47 -202
rect 75 -206 79 -202
rect 69 -213 73 -209
<< ndcontact >>
rect -6 -194 -2 -190
rect -6 -202 -2 -198
rect 33 -199 37 -195
rect 41 -199 45 -195
rect 53 -199 57 -195
rect 61 -199 65 -195
rect -6 -210 -2 -206
<< pdcontact >>
rect 33 -213 37 -209
rect 41 -213 45 -209
rect 53 -213 57 -209
rect 61 -213 65 -209
<< m2contact >>
rect 28 -180 32 -176
rect 48 -180 52 -176
rect -6 -187 -2 -183
rect 18 -196 22 -192
rect 61 -194 65 -190
rect 101 -194 105 -190
rect 28 -199 32 -195
rect 48 -199 52 -195
rect 18 -210 22 -206
<< psubstratepcontact >>
rect 34 -180 46 -176
<< nsubstratencontact >>
rect 79 -220 91 -216
use addsub  addsub_0
timestamp 1428972937
transform 1 0 58 0 1 -66
box -107 -58 97 79
<< end >>
