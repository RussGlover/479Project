magic
tech scmos
timestamp 1428277303
<< pwell >>
rect -78 8 -42 23
rect -25 8 0 25
rect -78 6 -46 8
<< nwell >>
rect -73 40 -63 43
rect -73 39 -50 40
rect -73 29 -10 39
<< polysilicon >>
rect -82 47 3 49
rect -82 42 -72 44
rect -65 36 -63 47
rect -48 42 3 44
rect -23 38 -21 42
rect -15 38 -13 40
rect -57 36 -55 38
rect -82 25 -71 27
rect -82 6 -80 8
rect -73 2 -71 25
rect -65 25 -63 32
rect -57 29 -55 32
rect -57 27 -47 29
rect -65 23 -55 25
rect -65 16 -63 18
rect -57 16 -55 23
rect -65 9 -63 12
rect -57 10 -55 12
rect -49 8 -47 27
rect -23 27 -21 34
rect -15 31 -13 34
rect -15 29 -5 31
rect -7 28 -5 29
rect -23 25 -13 27
rect -23 18 -21 20
rect -15 18 -13 25
rect -7 26 3 28
rect -23 13 -21 14
rect -62 6 -47 8
rect -41 11 -21 13
rect -15 12 -13 14
rect -41 2 -39 11
rect -23 10 -21 11
rect -7 10 -5 26
rect -23 8 -5 10
rect -7 6 3 8
rect -73 0 -39 2
<< ndiffusion >>
rect -66 12 -65 16
rect -63 12 -62 16
rect -58 12 -57 16
rect -55 12 -54 16
rect -24 14 -23 18
rect -21 14 -20 18
rect -16 14 -15 18
rect -13 14 -12 18
<< pdiffusion >>
rect -66 32 -65 36
rect -63 32 -62 36
rect -58 32 -57 36
rect -55 32 -54 36
rect -24 34 -23 38
rect -21 34 -20 38
rect -16 34 -15 38
rect -13 34 -12 38
<< metal1 >>
rect -68 40 -52 44
rect -74 32 -70 36
rect -50 32 -46 36
rect -32 34 -28 38
rect -8 34 -4 38
rect -20 33 -16 34
rect -62 31 -58 32
rect -50 22 -36 26
rect -20 18 -16 19
rect -62 16 -58 17
rect -74 12 -70 16
rect -50 12 -46 16
rect -32 14 -28 18
rect -8 14 -4 18
rect -20 10 -16 14
rect -78 8 -66 9
rect -76 5 -66 8
rect -34 6 -16 10
<< metal2 >>
rect -78 36 -74 50
rect -56 46 -52 50
rect -56 42 -42 46
rect -78 16 -74 32
rect -46 36 -42 42
rect -62 26 -58 27
rect -62 22 -54 26
rect -62 21 -58 22
rect -62 16 -58 17
rect -46 16 -42 32
rect -36 38 -32 39
rect -4 38 0 50
rect -36 26 -32 34
rect -36 18 -32 22
rect -20 33 -16 34
rect -20 23 -16 29
rect -20 18 -16 19
rect -4 18 0 34
rect -38 0 -34 6
<< ntransistor >>
rect -65 12 -63 16
rect -57 12 -55 16
rect -23 14 -21 18
rect -15 14 -13 18
<< ptransistor >>
rect -65 32 -63 36
rect -57 32 -55 36
rect -23 34 -21 38
rect -15 34 -13 38
<< polycontact >>
rect -72 40 -68 44
rect -52 40 -48 44
rect -80 4 -76 8
rect -66 5 -62 9
<< ndcontact >>
rect -70 12 -66 16
rect -62 12 -58 16
rect -54 12 -50 16
rect -28 14 -24 18
rect -20 14 -16 18
rect -12 14 -8 18
<< pdcontact >>
rect -70 32 -66 36
rect -62 32 -58 36
rect -54 32 -50 36
rect -28 34 -24 38
rect -20 34 -16 38
rect -12 34 -8 38
<< m2contact >>
rect -78 32 -74 36
rect -46 32 -42 36
rect -36 34 -32 38
rect -4 34 0 38
rect -62 27 -58 31
rect -20 29 -16 33
rect -54 22 -50 26
rect -36 22 -32 26
rect -62 17 -58 21
rect -20 19 -16 23
rect -78 12 -74 16
rect -46 12 -42 16
rect -36 14 -32 18
rect -4 14 0 18
rect -38 6 -34 10
<< psubstratepcontact >>
rect -78 19 -74 23
rect -4 21 0 25
<< end >>
