magic
tech scmos
timestamp 1428729313
<< pwell >>
rect -90 33 -77 46
rect -94 9 -78 33
<< nwell >>
rect -73 9 -57 46
<< polysilicon >>
rect -96 48 -75 49
rect -96 47 -79 48
rect -88 39 -86 41
rect -82 39 -72 41
rect -64 39 -62 41
rect -77 33 -75 39
rect -88 23 -86 25
rect -82 23 -69 25
rect -65 23 -57 25
rect -88 15 -86 17
rect -82 15 -69 17
rect -65 15 -57 17
<< ndiffusion >>
rect -86 41 -82 42
rect -86 38 -82 39
rect -86 25 -82 26
rect -86 17 -82 23
rect -86 14 -82 15
rect -86 9 -82 10
<< pdiffusion >>
rect -68 42 -64 46
rect -72 41 -64 42
rect -72 38 -64 39
rect -72 34 -68 38
rect -69 25 -65 26
rect -69 22 -65 23
rect -69 17 -65 18
rect -69 14 -65 15
rect -69 9 -65 10
<< metal1 >>
rect -94 38 -90 46
rect -82 44 -79 46
rect -75 44 -72 46
rect -82 42 -72 44
rect -61 38 -57 46
rect -94 34 -86 38
rect -64 34 -57 38
rect -94 22 -90 34
rect -82 29 -78 30
rect -74 29 -73 33
rect -61 30 -57 34
rect -82 26 -73 29
rect -65 26 -57 30
rect -78 22 -73 26
rect -61 22 -57 26
rect -73 18 -69 22
rect -94 14 -90 18
rect -61 14 -57 18
rect -94 10 -86 14
rect -65 10 -57 14
rect -94 9 -90 10
rect -61 9 -57 10
<< ntransistor >>
rect -86 39 -82 41
rect -86 23 -82 25
rect -86 15 -82 17
<< ptransistor >>
rect -72 39 -64 41
rect -69 23 -65 25
rect -69 15 -65 17
<< polycontact >>
rect -79 44 -75 48
rect -78 29 -74 33
<< ndcontact >>
rect -86 42 -82 46
rect -86 34 -82 38
rect -86 26 -82 30
rect -86 10 -82 14
<< pdcontact >>
rect -72 42 -68 46
rect -68 34 -64 38
rect -69 26 -65 30
rect -69 18 -65 22
rect -69 10 -65 14
<< m2contact >>
rect -78 18 -73 22
<< psubstratepcontact >>
rect -94 18 -90 22
<< nsubstratencontact >>
rect -61 18 -57 22
<< labels >>
rlabel polysilicon -96 47 -79 49 5 out
rlabel metal1 -94 22 -90 46 3 Gnd
rlabel metal1 -61 22 -57 46 7 Vdd
rlabel polysilicon -65 23 -57 25 7 A
rlabel polysilicon -65 15 -57 17 7 B
<< end >>
