magic
tech scmos
timestamp 1428739103
<< pwell >>
rect -89 54 -79 59
rect -89 41 -72 54
rect -89 9 -73 41
rect -89 7 -79 9
<< nwell >>
rect -68 9 -52 54
<< polysilicon >>
rect -91 56 -70 57
rect -91 55 -74 56
rect -83 47 -81 49
rect -77 47 -67 49
rect -59 47 -57 49
rect -72 41 -70 47
rect -83 31 -81 33
rect -77 31 -64 33
rect -60 31 -52 33
rect -83 23 -81 25
rect -77 23 -64 25
rect -60 23 -52 25
rect -83 15 -81 17
rect -77 15 -64 17
rect -60 15 -52 17
<< ndiffusion >>
rect -81 49 -77 50
rect -81 46 -77 47
rect -81 33 -77 34
rect -81 25 -77 31
rect -81 17 -77 23
rect -81 14 -77 15
rect -81 9 -77 10
<< pdiffusion >>
rect -63 50 -59 54
rect -67 49 -59 50
rect -67 46 -59 47
rect -67 42 -63 46
rect -64 33 -60 34
rect -64 30 -60 31
rect -64 25 -60 26
rect -64 22 -60 23
rect -64 17 -60 18
rect -64 14 -60 15
<< metal1 >>
rect -89 46 -85 54
rect -77 52 -74 54
rect -70 52 -67 54
rect -77 50 -67 52
rect -56 46 -52 54
rect -89 42 -81 46
rect -59 42 -52 46
rect -89 22 -85 42
rect -77 37 -73 38
rect -69 38 -68 41
rect -69 37 -64 38
rect -77 34 -64 37
rect -73 22 -68 34
rect -56 30 -52 42
rect -60 26 -52 30
rect -56 22 -52 26
rect -68 18 -64 22
rect -89 14 -85 18
rect -56 14 -52 18
rect -89 10 -81 14
rect -60 10 -52 14
rect -89 9 -85 10
rect -56 9 -52 10
<< ntransistor >>
rect -81 47 -77 49
rect -81 31 -77 33
rect -81 23 -77 25
rect -81 15 -77 17
<< ptransistor >>
rect -67 47 -59 49
rect -64 31 -60 33
rect -64 23 -60 25
rect -64 15 -60 17
<< polycontact >>
rect -74 52 -70 56
rect -73 37 -69 41
<< ndcontact >>
rect -81 50 -77 54
rect -81 42 -77 46
rect -81 34 -77 38
rect -81 10 -77 14
<< pdcontact >>
rect -67 50 -63 54
rect -63 42 -59 46
rect -64 34 -60 38
rect -64 26 -60 30
rect -64 18 -60 22
rect -64 10 -60 14
<< m2contact >>
rect -73 18 -68 22
<< psubstratepcontact >>
rect -89 18 -85 22
<< nsubstratencontact >>
rect -56 18 -52 22
<< labels >>
rlabel polysilicon -91 55 -74 57 5 out
rlabel polysilicon -83 31 -81 33 1 A
rlabel polysilicon -83 23 -81 25 1 B
rlabel polysilicon -83 15 -81 17 1 C
rlabel metal1 -89 22 -85 54 3 Gnd
rlabel metal1 -56 22 -52 54 7 Vdd
<< end >>
