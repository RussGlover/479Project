magic
tech scmos
timestamp 1428273030
<< nwell >>
rect -76 -24 88 20
<< polysilicon >>
rect -26 57 31 59
rect -65 49 -63 51
rect -37 49 -35 51
rect -26 49 -24 57
rect -22 53 21 55
rect -22 49 -20 53
rect -18 49 -16 51
rect -1 49 1 51
rect 8 49 10 51
rect 19 49 21 53
rect 29 49 31 57
rect 39 57 79 59
rect 39 49 41 57
rect 43 53 67 55
rect 43 49 45 53
rect 54 49 56 51
rect 65 49 67 53
rect 77 49 79 57
rect -65 17 -63 43
rect -65 -1 -63 13
rect -37 5 -35 43
rect -37 -1 -35 1
rect -26 -1 -24 43
rect -22 -1 -20 43
rect -18 19 -16 43
rect -1 26 1 43
rect 8 20 10 43
rect 19 37 21 43
rect 29 41 31 43
rect 39 41 41 43
rect 29 39 41 41
rect 43 37 45 43
rect 19 35 45 37
rect 40 34 44 35
rect 54 21 56 43
rect -18 17 8 19
rect -18 -1 -16 17
rect -1 -1 1 9
rect 8 -1 10 16
rect 19 5 45 7
rect 19 -1 21 5
rect 29 1 41 3
rect 29 -1 31 1
rect 39 -1 41 1
rect 43 -1 45 5
rect 54 -1 56 17
rect 65 -1 67 43
rect 77 41 79 43
rect 77 8 81 10
rect 77 -1 79 8
rect -65 -9 -63 -7
rect -37 -9 -35 -7
rect -26 -15 -24 -7
rect -22 -11 -20 -7
rect -18 -9 -16 -7
rect -1 -9 1 -7
rect 8 -9 10 -7
rect 19 -11 21 -7
rect -22 -13 21 -11
rect 29 -15 31 -7
rect -26 -17 31 -15
rect 39 -15 41 -7
rect 43 -11 45 -7
rect 54 -9 56 -7
rect 65 -11 67 -7
rect 43 -13 67 -11
rect 77 -15 79 -7
rect 39 -17 79 -15
<< ndiffusion >>
rect -76 48 -65 49
rect -76 43 -73 48
rect -69 43 -65 48
rect -63 48 -55 49
rect -63 44 -61 48
rect -57 44 -55 48
rect -63 43 -55 44
rect -49 48 -37 49
rect -49 44 -45 48
rect -41 44 -37 48
rect -49 43 -37 44
rect -35 48 -26 49
rect -35 44 -32 48
rect -28 44 -26 48
rect -35 43 -26 44
rect -24 43 -22 49
rect -20 43 -18 49
rect -16 48 -1 49
rect -16 44 -11 48
rect -7 44 -1 48
rect -16 43 -1 44
rect 1 48 8 49
rect 1 44 2 48
rect 6 44 8 48
rect 1 43 8 44
rect 10 48 19 49
rect 10 44 12 48
rect 16 44 19 48
rect 10 43 19 44
rect 21 48 29 49
rect 21 44 23 48
rect 27 44 29 48
rect 21 43 29 44
rect 31 48 39 49
rect 31 44 33 48
rect 37 44 39 48
rect 31 43 39 44
rect 41 43 43 49
rect 45 48 54 49
rect 45 44 47 48
rect 51 44 54 48
rect 45 43 54 44
rect 56 48 65 49
rect 56 44 58 48
rect 62 44 65 48
rect 56 43 65 44
rect 67 48 77 49
rect 67 44 69 48
rect 73 44 77 48
rect 67 43 77 44
rect 79 48 88 49
rect 79 44 82 48
rect 86 44 88 48
rect 79 43 88 44
<< pdiffusion >>
rect -76 -2 -65 -1
rect -76 -6 -73 -2
rect -69 -6 -65 -2
rect -76 -7 -65 -6
rect -63 -2 -55 -1
rect -63 -6 -61 -2
rect -57 -6 -55 -2
rect -63 -7 -55 -6
rect -49 -2 -37 -1
rect -49 -6 -45 -2
rect -41 -6 -37 -2
rect -49 -7 -37 -6
rect -35 -2 -26 -1
rect -35 -6 -32 -2
rect -28 -6 -26 -2
rect -35 -7 -26 -6
rect -24 -7 -22 -1
rect -20 -7 -18 -1
rect -16 -2 -1 -1
rect -16 -6 -11 -2
rect -7 -6 -1 -2
rect -16 -7 -1 -6
rect 1 -2 8 -1
rect 1 -6 2 -2
rect 6 -6 8 -2
rect 1 -7 8 -6
rect 10 -2 19 -1
rect 10 -6 12 -2
rect 16 -6 19 -2
rect 10 -7 19 -6
rect 21 -2 29 -1
rect 21 -6 23 -2
rect 27 -6 29 -2
rect 21 -7 29 -6
rect 31 -2 39 -1
rect 31 -6 33 -2
rect 37 -6 39 -2
rect 31 -7 39 -6
rect 41 -7 43 -1
rect 45 -2 54 -1
rect 45 -6 47 -2
rect 51 -6 54 -2
rect 45 -7 54 -6
rect 56 -2 65 -1
rect 56 -6 58 -2
rect 62 -6 65 -2
rect 56 -7 65 -6
rect 67 -2 77 -1
rect 67 -7 70 -2
rect 74 -7 77 -2
rect 79 -2 88 -1
rect 79 -6 82 -2
rect 86 -6 88 -2
rect 79 -7 88 -6
<< metal1 >>
rect -75 61 88 65
rect -61 48 -57 61
rect -32 48 -28 61
rect 12 48 16 61
rect 33 48 37 61
rect 69 48 73 61
rect -73 21 -69 44
rect -45 37 -41 44
rect -11 43 -7 44
rect 2 41 6 44
rect 23 41 27 44
rect 2 37 27 41
rect -4 33 40 34
rect -29 30 40 33
rect -29 29 -2 30
rect 47 27 51 44
rect 58 40 62 44
rect 82 40 86 44
rect 58 36 86 40
rect 3 24 51 27
rect 3 23 6 24
rect 3 22 5 23
rect -1 17 3 22
rect 47 20 52 21
rect -73 -2 -69 17
rect -62 13 3 17
rect 12 17 52 20
rect 56 17 78 21
rect 12 16 48 17
rect 3 9 51 13
rect 62 10 77 14
rect -45 -2 -41 5
rect -33 1 -11 5
rect -11 -2 -7 1
rect 2 1 27 5
rect 2 -2 6 1
rect 23 -2 27 1
rect 47 -2 51 9
rect 58 2 86 6
rect 58 -2 62 2
rect 82 -2 86 2
rect -61 -20 -57 -6
rect -32 -20 -28 -6
rect 12 -20 16 -6
rect 33 -20 37 -6
rect 70 -20 74 -6
rect -76 -24 88 -20
<< metal2 >>
rect -78 17 -73 21
rect -45 9 -41 33
rect -33 33 -29 71
rect -45 -33 -41 5
rect -22 -32 -18 71
rect -11 40 -7 43
rect -11 5 -7 36
rect -1 9 3 13
rect 30 -28 34 69
rect 58 14 62 71
rect 82 17 91 21
<< ntransistor >>
rect -65 43 -63 49
rect -37 43 -35 49
rect -26 43 -24 49
rect -22 43 -20 49
rect -18 43 -16 49
rect -1 43 1 49
rect 8 43 10 49
rect 19 43 21 49
rect 29 43 31 49
rect 39 43 41 49
rect 43 43 45 49
rect 54 43 56 49
rect 65 43 67 49
rect 77 43 79 49
<< ptransistor >>
rect -65 -7 -63 -1
rect -37 -7 -35 -1
rect -26 -7 -24 -1
rect -22 -7 -20 -1
rect -18 -7 -16 -1
rect -1 -7 1 -1
rect 8 -7 10 -1
rect 19 -7 21 -1
rect 29 -7 31 -1
rect 39 -7 41 -1
rect 43 -7 45 -1
rect 54 -7 56 -1
rect 65 -7 67 -1
rect 77 -7 79 -1
<< polycontact >>
rect -66 13 -62 17
rect -37 1 -33 5
rect -1 22 3 26
rect 40 30 44 34
rect 8 16 12 20
rect 52 17 56 21
rect -1 9 3 13
rect 77 10 81 14
<< ndcontact >>
rect -73 44 -69 48
rect -61 44 -57 48
rect -45 44 -41 48
rect -32 44 -28 48
rect -11 44 -7 48
rect 2 44 6 48
rect 12 44 16 48
rect 23 44 27 48
rect 33 44 37 48
rect 47 44 51 48
rect 58 44 62 48
rect 69 44 73 48
rect 82 44 86 48
<< pdcontact >>
rect -73 -6 -69 -2
rect -61 -6 -57 -2
rect -45 -6 -41 -2
rect -32 -6 -28 -2
rect -11 -6 -7 -2
rect 2 -6 6 -2
rect 12 -6 16 -2
rect 23 -6 27 -2
rect 33 -6 37 -2
rect 47 -6 51 -2
rect 58 -6 62 -2
rect 70 -6 74 -2
rect 82 -6 86 -2
<< m2contact >>
rect -45 33 -41 37
rect -11 36 -7 40
rect -33 29 -29 33
rect -73 17 -69 21
rect 78 17 82 21
rect 58 10 62 14
rect -45 5 -41 9
rect -11 1 -7 5
<< labels >>
rlabel metal2 -45 -33 -41 -33 1 Z
rlabel metal2 -78 17 -78 21 3 x
rlabel metal2 91 17 91 21 7 C
rlabel metal2 -33 71 -29 71 5 B
rlabel metal2 -22 -32 -18 -32 1 divideIn
rlabel metal2 30 69 34 69 5 fromShift
<< end >>
