magic
tech scmos
timestamp 1428802844
<< pwell >>
rect -74 286 -61 291
rect -74 276 -58 286
rect -80 272 -58 276
rect -87 259 -58 272
rect -85 244 -58 259
rect -87 231 -58 244
rect -85 218 -58 231
rect -87 215 -58 218
rect -87 205 -61 215
rect -74 190 -61 205
rect -87 178 -61 190
rect -87 177 -58 178
rect -74 168 -58 177
rect -88 165 -58 168
rect -88 132 -61 165
rect -74 125 -61 132
<< nwell >>
rect -107 258 -91 272
rect -53 265 -37 279
rect -107 231 -91 244
rect -52 227 -37 228
rect -107 204 -91 218
rect -53 215 -37 227
rect -107 168 -91 190
rect -107 137 -92 168
rect -53 165 -37 178
<< polysilicon >>
rect -89 320 -75 322
rect -89 266 -87 320
rect -37 296 -1 298
rect -37 288 7 290
rect -37 280 15 282
rect -102 264 -100 266
rect -92 264 -82 266
rect -78 264 -76 266
rect -104 260 -101 262
rect -103 258 -101 260
rect -103 256 -89 258
rect -104 252 -100 254
rect -102 248 -100 252
rect -102 246 -89 248
rect -73 241 -71 272
rect -37 246 -33 248
rect -76 240 -71 241
rect -77 239 -71 240
rect -102 237 -100 239
rect -92 237 -82 239
rect -78 238 -74 239
rect -37 238 -25 240
rect -78 237 -75 238
rect -37 230 -17 232
rect -144 228 -143 230
rect -89 220 -76 222
rect -89 212 -87 220
rect -102 210 -100 212
rect -92 210 -82 212
rect -78 210 -76 212
rect -104 206 -101 208
rect -103 204 -101 206
rect -103 202 -89 204
rect -104 198 -100 200
rect -102 194 -100 198
rect -37 196 -1 198
rect -102 192 -89 194
rect -37 188 7 190
rect -102 183 -100 185
rect -92 183 -82 185
rect -78 183 -76 185
rect -89 179 -87 183
rect -89 177 -83 179
rect -37 180 -9 182
rect -85 172 -83 177
rect -85 170 -73 172
rect -110 160 -101 162
rect -93 160 -83 162
rect -79 160 -77 162
rect -37 146 -17 148
rect -123 142 -101 144
rect -93 142 -83 144
rect -79 142 -77 144
rect -37 138 -25 140
rect -37 130 -33 132
<< ndiffusion >>
rect -82 266 -78 267
rect -82 263 -78 264
rect -82 239 -78 240
rect -82 236 -78 237
rect -82 212 -78 213
rect -82 209 -78 210
rect -82 185 -78 186
rect -82 182 -78 183
rect -83 162 -79 163
rect -83 159 -79 160
rect -83 144 -79 145
rect -83 141 -79 142
<< pdiffusion >>
rect -96 267 -92 271
rect -100 266 -92 267
rect -100 263 -92 264
rect -100 259 -96 263
rect -100 240 -96 244
rect -100 239 -92 240
rect -100 236 -92 237
rect -96 232 -92 236
rect -96 213 -92 217
rect -100 212 -92 213
rect -100 209 -92 210
rect -100 205 -96 209
rect -100 186 -96 190
rect -100 185 -92 186
rect -100 182 -92 183
rect -96 178 -92 182
rect -97 163 -93 167
rect -101 162 -93 163
rect -101 159 -93 160
rect -101 155 -97 159
rect -97 145 -93 149
rect -101 144 -93 145
rect -101 141 -93 142
rect -101 137 -97 141
<< metal1 >>
rect -455 328 -451 332
rect -246 314 -242 321
rect -234 307 -148 311
rect -325 300 -156 304
rect -164 292 -160 296
rect -455 288 -451 292
rect -164 285 -160 289
rect -164 278 -160 282
rect -107 271 -103 272
rect -74 271 -70 324
rect -107 267 -100 271
rect -78 267 -70 271
rect -455 229 -451 233
rect -148 231 -144 236
rect -141 212 -137 267
rect -107 236 -103 267
rect -92 259 -82 263
rect -89 258 -85 259
rect -89 244 -85 245
rect -92 240 -82 244
rect -74 236 -70 267
rect -107 232 -100 236
rect -78 232 -70 236
rect -107 217 -103 232
rect -74 217 -70 232
rect -107 213 -100 217
rect -78 213 -70 217
rect -455 189 -451 193
rect -107 182 -103 213
rect -92 205 -82 209
rect -89 204 -85 205
rect -89 190 -85 191
rect -92 186 -82 190
rect -74 182 -70 213
rect -107 178 -100 182
rect -78 178 -70 182
rect -152 170 -143 174
rect -107 167 -103 178
rect -74 167 -70 178
rect -117 160 -114 164
rect -107 163 -101 167
rect -79 163 -70 167
rect -455 149 -451 153
rect -164 152 -160 156
rect -107 149 -103 163
rect -93 155 -83 159
rect -90 150 -86 155
rect -74 149 -70 163
rect -199 132 -195 144
rect -455 128 -451 132
rect -327 128 -195 132
rect -157 118 -153 144
rect -127 140 -123 142
rect -107 145 -101 149
rect -79 145 -70 149
rect -107 139 -103 145
rect -93 137 -83 141
rect -90 136 -86 137
rect -90 130 -86 132
rect -90 126 -79 130
rect -98 110 -94 122
rect -83 98 -79 126
rect -74 120 -70 145
rect -41 121 -37 325
rect -33 250 -29 314
rect -33 134 -29 246
rect -25 142 -21 238
rect -25 102 -21 138
rect -17 150 -13 230
rect -9 184 -5 318
rect -1 207 3 296
rect -1 200 3 203
rect 7 192 11 288
rect 15 284 19 321
rect -17 110 -13 146
rect 7 122 11 188
rect 6 121 11 122
rect 6 94 10 121
<< metal2 >>
rect -156 174 -152 300
rect -148 240 -144 307
rect -157 160 -121 164
rect -117 160 -116 164
rect -290 140 -286 152
rect -199 148 -195 152
rect -157 148 -153 160
rect -195 144 -157 148
rect -290 136 -127 140
rect -345 128 -331 132
rect -290 121 -286 136
rect -338 116 -286 121
rect -166 94 -162 136
rect -90 126 -86 154
rect -94 122 -86 126
rect -1 118 3 203
rect -153 114 3 118
rect -94 106 -17 110
rect -83 98 -25 102
rect -166 90 6 94
<< ntransistor >>
rect -82 264 -78 266
rect -82 237 -78 239
rect -82 210 -78 212
rect -82 183 -78 185
rect -83 160 -79 162
rect -83 142 -79 144
<< ptransistor >>
rect -100 264 -92 266
rect -100 237 -92 239
rect -100 210 -92 212
rect -100 183 -92 185
rect -101 160 -93 162
rect -101 142 -93 144
<< polycontact >>
rect -1 296 3 300
rect 7 288 11 292
rect 15 280 19 284
rect -89 254 -85 258
rect -89 245 -85 249
rect -33 246 -29 250
rect -25 238 -21 242
rect -148 227 -144 231
rect -17 230 -13 234
rect -89 200 -85 204
rect -1 196 3 200
rect -89 191 -85 195
rect 7 188 11 192
rect -9 180 -5 184
rect -143 170 -139 174
rect -114 160 -110 164
rect -127 142 -123 146
rect -17 146 -13 150
rect -25 138 -21 142
rect -90 132 -86 136
rect -33 130 -29 134
<< ndcontact >>
rect -82 267 -78 271
rect -82 259 -78 263
rect -82 240 -78 244
rect -82 232 -78 236
rect -82 213 -78 217
rect -82 205 -78 209
rect -82 186 -78 190
rect -82 178 -78 182
rect -83 163 -79 167
rect -83 155 -79 159
rect -83 145 -79 149
rect -83 137 -79 141
<< pdcontact >>
rect -100 267 -96 271
rect -96 259 -92 263
rect -96 240 -92 244
rect -100 232 -96 236
rect -100 213 -96 217
rect -96 205 -92 209
rect -96 186 -92 190
rect -100 178 -96 182
rect -101 163 -97 167
rect -97 155 -93 159
rect -101 145 -97 149
rect -97 137 -93 141
<< m2contact >>
rect -238 307 -234 311
rect -148 307 -144 311
rect -329 300 -325 304
rect -156 300 -152 304
rect -148 236 -144 240
rect -156 170 -152 174
rect -121 160 -117 164
rect -199 144 -195 148
rect -349 128 -345 132
rect -331 128 -327 132
rect -157 144 -153 148
rect -342 116 -338 121
rect -127 136 -123 140
rect -157 114 -153 118
rect -98 122 -94 126
rect -98 106 -94 110
rect -1 203 3 207
rect -17 106 -13 110
rect -25 98 -21 102
rect 6 90 10 94
use controller_part2  controller_part2_0
timestamp 1428732039
transform 1 0 -331 0 1 283
box -120 -190 -7 50
use reg2bit2  reg2bit2_0
timestamp 1428802636
transform 1 0 -316 0 1 310
box -17 -158 156 8
use and3gate  and3gate_3
timestamp 1428739103
transform 1 0 15 0 1 265
box -91 7 -52 59
use andgate  andgate_1
timestamp 1428729313
transform 1 0 -47 0 -1 277
box -96 9 -57 49
use and3gate  and3gate_0
timestamp 1428739103
transform 1 0 15 0 1 215
box -91 7 -52 59
use andgate  andgate_0
timestamp 1428729313
transform 1 0 -47 0 -1 223
box -96 9 -57 49
use and3gate  and3gate_1
timestamp 1428739103
transform 1 0 15 0 1 165
box -91 7 -52 59
use and3gate  and3gate_2
timestamp 1428739103
transform 1 0 15 0 1 115
box -91 7 -52 59
<< labels >>
rlabel metal1 7 192 11 288 7 B
rlabel metal1 -17 150 -13 198 1 An
rlabel metal1 -25 142 -21 198 1 Bn
rlabel metal1 -33 134 -29 198 1 Startn
rlabel metal1 -147 170 -143 174 3 Bout
rlabel metal1 -74 287 -70 324 1 Gnd
rlabel metal1 -41 319 -37 324 5 Vdd
rlabel metal1 -141 214 -137 267 1 Gnd
rlabel metal1 -1 200 3 296 1 A
rlabel metal1 -9 184 -5 280 1 Signn
rlabel metal1 -107 177 -103 272 1 Vdd2
rlabel metal1 15 284 19 321 7 sign
rlabel metal1 -148 231 -144 236 1 Aout
rlabel metal1 -455 128 -451 132 3 inbit
rlabel metal1 -455 149 -451 153 3 shift
rlabel metal1 -455 189 -451 193 3 sel0
rlabel metal1 -455 229 -451 233 3 s1
rlabel metal1 -455 288 -451 292 3 add
rlabel metal1 -455 328 -451 332 4 load
rlabel metal1 -246 314 -242 321 1 Vdd
rlabel metal1 -164 278 -160 282 1 rst
rlabel metal1 -164 285 -160 289 1 Clkn
rlabel metal1 -164 292 -160 296 1 Clk
rlabel metal1 -164 152 -160 156 1 Gnd
<< end >>
