magic
tech scmos
timestamp 1428304724
<< pwell >>
rect 24 -111 126 -71
rect 193 -111 295 -71
rect 24 -119 48 -111
rect 193 -119 217 -111
<< nwell >>
rect 73 -131 126 -115
rect 242 -131 295 -115
<< polysilicon >>
rect 12 -98 28 -96
rect 32 -98 60 -96
rect 181 -98 197 -96
rect 201 -98 229 -96
rect 86 -103 88 -101
rect 110 -103 112 -101
rect 255 -103 257 -101
rect 279 -103 281 -101
rect 20 -106 28 -104
rect 32 -106 68 -104
rect 189 -106 197 -104
rect 201 -106 237 -104
rect 86 -111 88 -107
rect 110 -111 112 -107
rect 255 -111 257 -107
rect 279 -111 281 -107
rect 86 -119 88 -115
rect 110 -119 112 -115
rect 255 -119 257 -115
rect 279 -119 281 -115
rect 86 -125 88 -123
rect 110 -125 112 -123
rect 255 -125 257 -123
rect 279 -125 281 -123
<< ndiffusion >>
rect 28 -96 32 -95
rect 28 -99 32 -98
rect 197 -96 201 -95
rect 197 -99 201 -98
rect 28 -104 32 -103
rect 28 -107 32 -106
rect 85 -107 86 -103
rect 88 -107 89 -103
rect 109 -107 110 -103
rect 112 -107 113 -103
rect 197 -104 201 -103
rect 197 -107 201 -106
rect 254 -107 255 -103
rect 257 -107 258 -103
rect 278 -107 279 -103
rect 281 -107 282 -103
<< pdiffusion >>
rect 85 -123 86 -119
rect 88 -123 89 -119
rect 109 -123 110 -119
rect 112 -123 113 -119
rect 254 -123 255 -119
rect 257 -123 258 -119
rect 278 -123 279 -119
rect 281 -123 282 -119
<< metal1 >>
rect -18 -77 76 -73
rect 80 -77 84 -73
rect 96 -77 100 -73
rect 104 -77 245 -73
rect 249 -77 253 -73
rect 265 -77 269 -73
rect 273 -77 315 -73
rect -18 -85 28 -81
rect 40 -85 197 -81
rect 209 -85 315 -81
rect -18 -92 12 -88
rect 8 -95 12 -92
rect 28 -91 32 -85
rect 60 -92 181 -88
rect 60 -95 64 -92
rect 177 -95 181 -92
rect 197 -91 201 -85
rect 229 -92 315 -88
rect 229 -95 233 -92
rect -18 -99 -2 -95
rect 68 -99 167 -95
rect 237 -99 315 -95
rect -6 -111 -2 -99
rect 32 -103 48 -99
rect 16 -111 20 -107
rect 32 -111 36 -107
rect 44 -111 48 -103
rect 68 -103 72 -99
rect 80 -107 81 -103
rect 93 -111 97 -103
rect 104 -107 105 -103
rect 117 -111 121 -103
rect 163 -111 167 -99
rect 201 -103 217 -99
rect 185 -111 189 -107
rect 201 -111 205 -107
rect 213 -111 217 -103
rect 237 -103 241 -99
rect 249 -107 250 -103
rect 262 -111 266 -103
rect 273 -107 274 -103
rect 286 -111 290 -103
rect -6 -115 20 -111
rect 44 -115 85 -111
rect 93 -115 109 -111
rect 117 -115 122 -111
rect 163 -115 189 -111
rect 213 -115 254 -111
rect 262 -115 278 -111
rect 286 -115 291 -111
rect 93 -123 97 -115
rect 117 -123 121 -115
rect 262 -123 266 -115
rect 286 -123 290 -115
rect 81 -127 85 -123
rect 105 -127 109 -123
rect 250 -127 254 -123
rect 274 -127 278 -123
rect -18 -131 89 -127
rect 101 -131 258 -127
rect 270 -131 315 -127
<< metal2 >>
rect 28 -81 32 -73
rect 36 -107 40 -85
rect 76 -103 80 -77
rect 100 -103 104 -77
rect 122 -111 126 -73
rect 197 -81 201 -73
rect 205 -107 209 -85
rect 245 -103 249 -77
rect 269 -103 273 -77
rect 291 -111 295 -73
<< ntransistor >>
rect 28 -98 32 -96
rect 197 -98 201 -96
rect 28 -106 32 -104
rect 86 -107 88 -103
rect 110 -107 112 -103
rect 197 -106 201 -104
rect 255 -107 257 -103
rect 279 -107 281 -103
<< ptransistor >>
rect 86 -123 88 -119
rect 110 -123 112 -119
rect 255 -123 257 -119
rect 279 -123 281 -119
<< polycontact >>
rect 8 -99 12 -95
rect 60 -99 64 -95
rect 177 -99 181 -95
rect 229 -99 233 -95
rect 16 -107 20 -103
rect 68 -107 72 -103
rect 185 -107 189 -103
rect 237 -107 241 -103
rect 85 -115 89 -111
rect 109 -115 113 -111
rect 254 -115 258 -111
rect 278 -115 282 -111
<< ndcontact >>
rect 28 -95 32 -91
rect 197 -95 201 -91
rect 28 -103 32 -99
rect 197 -103 201 -99
rect 81 -107 85 -103
rect 89 -107 93 -103
rect 105 -107 109 -103
rect 113 -107 117 -103
rect 250 -107 254 -103
rect 258 -107 262 -103
rect 274 -107 278 -103
rect 282 -107 286 -103
rect 28 -111 32 -107
rect 197 -111 201 -107
<< pdcontact >>
rect 81 -123 85 -119
rect 89 -123 93 -119
rect 105 -123 109 -119
rect 113 -123 117 -119
rect 250 -123 254 -119
rect 258 -123 262 -119
rect 274 -123 278 -119
rect 282 -123 286 -119
<< m2contact >>
rect 76 -77 80 -73
rect 100 -77 104 -73
rect 245 -77 249 -73
rect 269 -77 273 -73
rect 28 -85 32 -81
rect 36 -85 40 -81
rect 197 -85 201 -81
rect 205 -85 209 -81
rect 36 -111 40 -107
rect 76 -107 80 -103
rect 100 -107 104 -103
rect 205 -111 209 -107
rect 245 -107 249 -103
rect 269 -107 273 -103
rect 122 -115 126 -111
rect 291 -115 295 -111
<< psubstratepcontact >>
rect 84 -77 96 -73
rect 253 -77 265 -73
<< nsubstratencontact >>
rect 89 -131 101 -127
rect 258 -131 270 -127
<< labels >>
rlabel metal1 313 -75 313 -75 6 GND
rlabel metal1 313 -129 313 -129 8 Vdd
rlabel metal2 293 -75 293 -75 5 OUT0
rlabel metal1 313 -90 313 -90 7 ShiftB
rlabel metal1 313 -97 313 -97 7 Shift
rlabel metal2 124 -75 124 -75 5 OUT1
rlabel metal2 199 -75 199 -75 5 IN1
rlabel metal1 313 -83 313 -83 7 IN0
rlabel metal2 30 -75 30 -75 5 IN2
<< end >>
