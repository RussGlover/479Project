magic
tech scmos
timestamp 1428732039
<< pwell >>
rect -101 33 -72 50
rect -101 10 -73 33
rect -101 -7 -72 10
rect -101 -30 -73 -7
rect -101 -47 -72 -30
rect -101 -70 -73 -47
rect -101 -87 -72 -70
rect -101 -110 -73 -87
rect -101 -127 -72 -110
rect -101 -150 -73 -127
rect -101 -167 -72 -150
rect -101 -190 -73 -167
rect -38 -190 -22 50
<< nwell >>
rect -119 -190 -104 50
rect -68 -190 -40 50
<< polysilicon >>
rect -92 48 -70 49
rect -92 47 -74 48
rect -83 39 -81 41
rect -77 39 -67 41
rect -59 39 -57 41
rect -51 39 -48 41
rect -44 39 -34 41
rect -30 39 -18 41
rect -72 33 -70 39
rect -54 31 -41 33
rect -54 25 -52 31
rect -89 23 -81 25
rect -77 23 -64 25
rect -60 23 -52 25
rect -50 19 -48 21
rect -44 19 -34 21
rect -30 19 -11 21
rect -89 15 -81 17
rect -77 15 -64 17
rect -60 15 -52 17
rect -54 13 -52 15
rect -54 11 -41 13
rect -92 8 -70 9
rect -92 7 -74 8
rect -83 -1 -81 1
rect -77 -1 -67 1
rect -59 -1 -57 1
rect -51 -1 -48 1
rect -44 -1 -34 1
rect -30 -1 -18 1
rect -72 -7 -70 -1
rect -54 -9 -41 -7
rect -54 -15 -52 -9
rect -89 -17 -81 -15
rect -77 -17 -64 -15
rect -60 -17 -52 -15
rect -43 -21 -11 -19
rect -89 -25 -81 -23
rect -77 -25 -64 -23
rect -60 -25 -52 -23
rect -54 -27 -52 -25
rect -43 -27 -41 -21
rect -54 -29 -41 -27
rect -103 -32 -70 -31
rect -103 -33 -74 -32
rect -103 -39 -101 -33
rect -113 -41 -111 -39
rect -107 -41 -96 -39
rect -92 -41 -90 -39
rect -83 -41 -81 -39
rect -77 -41 -67 -39
rect -59 -41 -57 -39
rect -51 -41 -48 -39
rect -44 -41 -34 -39
rect -30 -41 -18 -39
rect -72 -47 -70 -41
rect -54 -49 -41 -47
rect -54 -55 -52 -49
rect -89 -57 -81 -55
rect -77 -57 -64 -55
rect -60 -57 -52 -55
rect -50 -61 -48 -59
rect -44 -61 -34 -59
rect -30 -61 -11 -59
rect -89 -65 -81 -63
rect -77 -65 -64 -63
rect -60 -65 -52 -63
rect -54 -67 -52 -65
rect -54 -69 -41 -67
rect -103 -72 -70 -71
rect -103 -73 -74 -72
rect -103 -79 -101 -73
rect -113 -81 -111 -79
rect -107 -81 -96 -79
rect -92 -81 -90 -79
rect -83 -81 -81 -79
rect -77 -81 -67 -79
rect -59 -81 -57 -79
rect -32 -81 -18 -79
rect -72 -87 -70 -81
rect -32 -87 -30 -81
rect -54 -89 -30 -87
rect -54 -95 -52 -89
rect -89 -97 -81 -95
rect -77 -97 -64 -95
rect -60 -97 -52 -95
rect -50 -101 -48 -99
rect -44 -101 -34 -99
rect -30 -101 -11 -99
rect -89 -105 -81 -103
rect -77 -105 -64 -103
rect -60 -105 -52 -103
rect -54 -107 -52 -105
rect -54 -109 -41 -107
rect -103 -112 -70 -111
rect -103 -113 -74 -112
rect -103 -119 -101 -113
rect -113 -121 -111 -119
rect -107 -121 -96 -119
rect -92 -121 -90 -119
rect -83 -121 -81 -119
rect -77 -121 -67 -119
rect -59 -121 -57 -119
rect -32 -121 -18 -119
rect -72 -127 -70 -121
rect -32 -127 -30 -121
rect -54 -129 -30 -127
rect -54 -135 -52 -129
rect -89 -137 -81 -135
rect -77 -137 -64 -135
rect -60 -137 -52 -135
rect -32 -141 -11 -139
rect -89 -145 -81 -143
rect -77 -145 -64 -143
rect -60 -145 -52 -143
rect -54 -147 -52 -145
rect -32 -147 -30 -141
rect -54 -149 -30 -147
rect -92 -152 -70 -151
rect -92 -153 -74 -152
rect -83 -161 -81 -159
rect -77 -161 -67 -159
rect -59 -161 -57 -159
rect -32 -161 -18 -159
rect -72 -167 -70 -161
rect -32 -167 -30 -161
rect -54 -169 -30 -167
rect -54 -175 -52 -169
rect -89 -177 -81 -175
rect -77 -177 -64 -175
rect -60 -177 -52 -175
rect -50 -181 -48 -179
rect -44 -181 -34 -179
rect -30 -181 -11 -179
rect -89 -185 -81 -183
rect -77 -185 -64 -183
rect -60 -185 -52 -183
rect -54 -187 -52 -185
rect -54 -189 -41 -187
<< ndiffusion >>
rect -81 41 -77 42
rect -34 41 -30 42
rect -81 38 -77 39
rect -34 38 -30 39
rect -81 25 -77 26
rect -81 17 -77 23
rect -34 21 -30 22
rect -81 14 -77 15
rect -34 18 -30 19
rect -81 1 -77 2
rect -34 1 -30 2
rect -81 -2 -77 -1
rect -34 -2 -30 -1
rect -81 -15 -77 -14
rect -81 -23 -77 -17
rect -81 -26 -77 -25
rect -96 -39 -92 -38
rect -81 -39 -77 -38
rect -34 -39 -30 -38
rect -96 -42 -92 -41
rect -81 -42 -77 -41
rect -34 -42 -30 -41
rect -81 -55 -77 -54
rect -81 -63 -77 -57
rect -34 -59 -30 -58
rect -81 -66 -77 -65
rect -34 -62 -30 -61
rect -96 -79 -92 -78
rect -81 -79 -77 -78
rect -96 -82 -92 -81
rect -81 -82 -77 -81
rect -81 -95 -77 -94
rect -81 -103 -77 -97
rect -34 -99 -30 -98
rect -81 -106 -77 -105
rect -34 -102 -30 -101
rect -96 -119 -92 -118
rect -81 -119 -77 -118
rect -96 -122 -92 -121
rect -81 -122 -77 -121
rect -81 -135 -77 -134
rect -81 -143 -77 -137
rect -81 -146 -77 -145
rect -81 -159 -77 -158
rect -81 -162 -77 -161
rect -81 -175 -77 -174
rect -81 -183 -77 -177
rect -34 -179 -30 -178
rect -81 -186 -77 -185
rect -34 -182 -30 -181
<< pdiffusion >>
rect -63 42 -59 46
rect -67 41 -59 42
rect -48 41 -44 42
rect -67 38 -59 39
rect -67 34 -63 38
rect -48 38 -44 39
rect -64 25 -60 26
rect -64 22 -60 23
rect -48 21 -44 22
rect -48 18 -44 19
rect -64 17 -60 18
rect -64 14 -60 15
rect -63 2 -59 6
rect -67 1 -59 2
rect -48 1 -44 2
rect -67 -2 -59 -1
rect -67 -6 -63 -2
rect -48 -2 -44 -1
rect -64 -15 -60 -14
rect -64 -18 -60 -17
rect -64 -23 -60 -22
rect -64 -26 -60 -25
rect -111 -39 -107 -38
rect -63 -38 -59 -34
rect -67 -39 -59 -38
rect -48 -39 -44 -38
rect -111 -42 -107 -41
rect -67 -42 -59 -41
rect -67 -46 -63 -42
rect -48 -42 -44 -41
rect -64 -55 -60 -54
rect -64 -58 -60 -57
rect -48 -59 -44 -58
rect -48 -62 -44 -61
rect -64 -63 -60 -62
rect -64 -66 -60 -65
rect -111 -79 -107 -78
rect -63 -78 -59 -74
rect -67 -79 -59 -78
rect -111 -82 -107 -81
rect -67 -82 -59 -81
rect -67 -86 -63 -82
rect -64 -95 -60 -94
rect -64 -98 -60 -97
rect -48 -99 -44 -98
rect -48 -102 -44 -101
rect -64 -103 -60 -102
rect -64 -106 -60 -105
rect -111 -119 -107 -118
rect -63 -118 -59 -114
rect -67 -119 -59 -118
rect -111 -122 -107 -121
rect -67 -122 -59 -121
rect -67 -126 -63 -122
rect -64 -135 -60 -134
rect -64 -138 -60 -137
rect -64 -143 -60 -142
rect -64 -146 -60 -145
rect -63 -158 -59 -154
rect -67 -159 -59 -158
rect -67 -162 -59 -161
rect -67 -166 -63 -162
rect -64 -175 -60 -174
rect -64 -178 -60 -177
rect -48 -179 -44 -178
rect -48 -182 -44 -181
rect -64 -183 -60 -182
rect -64 -186 -60 -185
<< metal1 >>
rect -120 45 -96 49
rect -89 38 -85 50
rect -77 44 -74 46
rect -56 46 -52 50
rect -26 46 -22 50
rect -70 44 -67 46
rect -77 42 -67 44
rect -56 42 -48 46
rect -30 42 -22 46
rect -56 38 -52 42
rect -89 34 -81 38
rect -59 34 -52 38
rect -44 34 -34 38
rect -89 22 -85 34
rect -77 29 -73 30
rect -69 29 -68 33
rect -56 30 -52 34
rect -77 26 -68 29
rect -60 26 -52 30
rect -26 26 -22 42
rect -73 22 -68 26
rect -56 22 -48 26
rect -30 22 -22 26
rect -68 18 -64 22
rect -89 14 -85 18
rect -56 14 -52 18
rect -44 14 -34 18
rect -89 10 -81 14
rect -60 10 -52 14
rect -120 5 -96 9
rect -89 -2 -85 10
rect -77 4 -74 6
rect -56 6 -52 10
rect -26 6 -22 22
rect -70 4 -67 6
rect -77 2 -67 4
rect -56 2 -48 6
rect -30 2 -22 6
rect -56 -2 -52 2
rect -89 -6 -81 -2
rect -59 -6 -52 -2
rect -44 -6 -34 -2
rect -89 -18 -85 -6
rect -77 -11 -73 -10
rect -69 -11 -68 -7
rect -56 -10 -52 -6
rect -77 -14 -68 -11
rect -60 -14 -52 -10
rect -73 -18 -68 -14
rect -56 -18 -52 -14
rect -68 -22 -64 -18
rect -89 -26 -85 -22
rect -56 -26 -52 -22
rect -89 -30 -81 -26
rect -60 -30 -52 -26
rect -89 -34 -85 -30
rect -115 -38 -111 -34
rect -92 -38 -85 -34
rect -77 -36 -74 -34
rect -56 -34 -52 -30
rect -26 -34 -22 2
rect -70 -36 -67 -34
rect -77 -38 -67 -36
rect -56 -38 -48 -34
rect -30 -38 -22 -34
rect -89 -42 -85 -38
rect -56 -42 -52 -38
rect -107 -46 -96 -42
rect -89 -46 -81 -42
rect -59 -46 -52 -42
rect -44 -46 -34 -42
rect -104 -50 -100 -46
rect -120 -54 -100 -50
rect -89 -58 -85 -46
rect -77 -51 -73 -50
rect -69 -51 -68 -47
rect -56 -50 -52 -46
rect -77 -54 -68 -51
rect -60 -54 -52 -50
rect -26 -54 -22 -38
rect -73 -58 -68 -54
rect -56 -58 -48 -54
rect -30 -58 -22 -54
rect -68 -62 -64 -58
rect -89 -66 -85 -62
rect -56 -66 -52 -62
rect -44 -66 -34 -62
rect -89 -70 -81 -66
rect -60 -70 -52 -66
rect -89 -74 -85 -70
rect -115 -78 -111 -74
rect -92 -78 -85 -74
rect -77 -76 -74 -74
rect -70 -76 -67 -74
rect -77 -78 -67 -76
rect -89 -82 -85 -78
rect -56 -82 -52 -70
rect -107 -86 -96 -82
rect -89 -86 -81 -82
rect -59 -86 -52 -82
rect -104 -90 -100 -86
rect -120 -94 -100 -90
rect -89 -98 -85 -86
rect -77 -91 -73 -90
rect -69 -91 -68 -87
rect -56 -90 -52 -86
rect -77 -94 -68 -91
rect -60 -94 -52 -90
rect -26 -94 -22 -58
rect -73 -98 -68 -94
rect -56 -98 -48 -94
rect -30 -98 -22 -94
rect -68 -102 -64 -98
rect -89 -106 -85 -102
rect -56 -106 -52 -102
rect -44 -106 -34 -102
rect -89 -110 -81 -106
rect -60 -110 -52 -106
rect -89 -114 -85 -110
rect -115 -118 -111 -114
rect -92 -118 -85 -114
rect -77 -116 -74 -114
rect -70 -116 -67 -114
rect -77 -118 -67 -116
rect -89 -122 -85 -118
rect -56 -122 -52 -110
rect -107 -126 -96 -122
rect -89 -126 -81 -122
rect -59 -126 -52 -122
rect -104 -130 -100 -126
rect -120 -134 -100 -130
rect -89 -138 -85 -126
rect -77 -131 -73 -130
rect -69 -131 -68 -127
rect -56 -130 -52 -126
rect -77 -134 -68 -131
rect -60 -134 -52 -130
rect -73 -138 -68 -134
rect -56 -138 -52 -134
rect -68 -142 -64 -138
rect -89 -146 -85 -142
rect -56 -146 -52 -142
rect -89 -150 -81 -146
rect -60 -150 -52 -146
rect -120 -155 -96 -151
rect -89 -162 -85 -150
rect -77 -156 -74 -154
rect -70 -156 -67 -154
rect -77 -158 -67 -156
rect -56 -162 -52 -150
rect -89 -166 -81 -162
rect -59 -166 -52 -162
rect -119 -190 -115 -177
rect -89 -178 -85 -166
rect -77 -171 -73 -170
rect -69 -171 -68 -167
rect -56 -170 -52 -166
rect -77 -174 -68 -171
rect -60 -174 -52 -170
rect -26 -174 -22 -98
rect -73 -178 -68 -174
rect -56 -178 -48 -174
rect -30 -178 -22 -174
rect -68 -182 -64 -178
rect -89 -186 -85 -182
rect -56 -186 -52 -182
rect -44 -186 -34 -182
rect -89 -190 -81 -186
rect -60 -190 -52 -186
rect -26 -190 -22 -178
rect -18 42 -14 50
rect -18 2 -14 38
rect -18 -38 -14 -2
rect -18 -78 -14 -42
rect -18 -118 -14 -82
rect -18 -158 -14 -122
rect -18 -190 -14 -162
rect -11 22 -7 50
rect -11 -18 -7 18
rect -11 -58 -7 -22
rect -11 -98 -7 -62
rect -11 -138 -7 -102
rect -11 -178 -7 -142
rect -11 -190 -7 -182
<< metal2 >>
rect -119 -74 -115 -38
rect -119 -114 -115 -78
rect -119 -173 -115 -118
<< ntransistor >>
rect -81 39 -77 41
rect -34 39 -30 41
rect -81 23 -77 25
rect -34 19 -30 21
rect -81 15 -77 17
rect -81 -1 -77 1
rect -34 -1 -30 1
rect -81 -17 -77 -15
rect -81 -25 -77 -23
rect -96 -41 -92 -39
rect -81 -41 -77 -39
rect -34 -41 -30 -39
rect -81 -57 -77 -55
rect -34 -61 -30 -59
rect -81 -65 -77 -63
rect -96 -81 -92 -79
rect -81 -81 -77 -79
rect -81 -97 -77 -95
rect -34 -101 -30 -99
rect -81 -105 -77 -103
rect -96 -121 -92 -119
rect -81 -121 -77 -119
rect -81 -137 -77 -135
rect -81 -145 -77 -143
rect -81 -161 -77 -159
rect -81 -177 -77 -175
rect -34 -181 -30 -179
rect -81 -185 -77 -183
<< ptransistor >>
rect -67 39 -59 41
rect -48 39 -44 41
rect -64 23 -60 25
rect -48 19 -44 21
rect -64 15 -60 17
rect -67 -1 -59 1
rect -48 -1 -44 1
rect -64 -17 -60 -15
rect -64 -25 -60 -23
rect -111 -41 -107 -39
rect -67 -41 -59 -39
rect -48 -41 -44 -39
rect -64 -57 -60 -55
rect -48 -61 -44 -59
rect -64 -65 -60 -63
rect -111 -81 -107 -79
rect -67 -81 -59 -79
rect -64 -97 -60 -95
rect -48 -101 -44 -99
rect -64 -105 -60 -103
rect -111 -121 -107 -119
rect -67 -121 -59 -119
rect -64 -137 -60 -135
rect -64 -145 -60 -143
rect -67 -161 -59 -159
rect -64 -177 -60 -175
rect -48 -181 -44 -179
rect -64 -185 -60 -183
<< polycontact >>
rect -96 45 -92 49
rect -74 44 -70 48
rect -18 38 -14 42
rect -73 29 -69 33
rect -41 30 -37 34
rect -11 18 -7 22
rect -41 10 -37 14
rect -96 5 -92 9
rect -74 4 -70 8
rect -18 -2 -14 2
rect -73 -11 -69 -7
rect -41 -10 -37 -6
rect -11 -22 -7 -18
rect -74 -36 -70 -32
rect -18 -42 -14 -38
rect -73 -51 -69 -47
rect -41 -50 -37 -46
rect -11 -62 -7 -58
rect -41 -70 -37 -66
rect -74 -76 -70 -72
rect -18 -82 -14 -78
rect -73 -91 -69 -87
rect -11 -102 -7 -98
rect -41 -110 -37 -106
rect -74 -116 -70 -112
rect -18 -122 -14 -118
rect -73 -131 -69 -127
rect -11 -142 -7 -138
rect -96 -155 -92 -151
rect -74 -156 -70 -152
rect -18 -162 -14 -158
rect -73 -171 -69 -167
rect -11 -182 -7 -178
rect -41 -190 -37 -186
<< ndcontact >>
rect -81 42 -77 46
rect -34 42 -30 46
rect -81 34 -77 38
rect -34 34 -30 38
rect -81 26 -77 30
rect -34 22 -30 26
rect -81 10 -77 14
rect -34 14 -30 18
rect -81 2 -77 6
rect -34 2 -30 6
rect -81 -6 -77 -2
rect -34 -6 -30 -2
rect -81 -14 -77 -10
rect -81 -30 -77 -26
rect -96 -38 -92 -34
rect -81 -38 -77 -34
rect -34 -38 -30 -34
rect -96 -46 -92 -42
rect -81 -46 -77 -42
rect -34 -46 -30 -42
rect -81 -54 -77 -50
rect -34 -58 -30 -54
rect -81 -70 -77 -66
rect -34 -66 -30 -62
rect -96 -78 -92 -74
rect -81 -78 -77 -74
rect -96 -86 -92 -82
rect -81 -86 -77 -82
rect -81 -94 -77 -90
rect -34 -98 -30 -94
rect -81 -110 -77 -106
rect -34 -106 -30 -102
rect -96 -118 -92 -114
rect -81 -118 -77 -114
rect -96 -126 -92 -122
rect -81 -126 -77 -122
rect -81 -134 -77 -130
rect -81 -150 -77 -146
rect -81 -158 -77 -154
rect -81 -166 -77 -162
rect -81 -174 -77 -170
rect -34 -178 -30 -174
rect -81 -190 -77 -186
rect -34 -186 -30 -182
<< pdcontact >>
rect -67 42 -63 46
rect -48 42 -44 46
rect -63 34 -59 38
rect -48 34 -44 38
rect -64 26 -60 30
rect -48 22 -44 26
rect -64 18 -60 22
rect -64 10 -60 14
rect -48 14 -44 18
rect -67 2 -63 6
rect -48 2 -44 6
rect -63 -6 -59 -2
rect -48 -6 -44 -2
rect -64 -14 -60 -10
rect -64 -22 -60 -18
rect -64 -30 -60 -26
rect -111 -38 -107 -34
rect -67 -38 -63 -34
rect -48 -38 -44 -34
rect -111 -46 -107 -42
rect -63 -46 -59 -42
rect -48 -46 -44 -42
rect -64 -54 -60 -50
rect -48 -58 -44 -54
rect -64 -62 -60 -58
rect -64 -70 -60 -66
rect -48 -66 -44 -62
rect -111 -78 -107 -74
rect -67 -78 -63 -74
rect -111 -86 -107 -82
rect -63 -86 -59 -82
rect -64 -94 -60 -90
rect -48 -98 -44 -94
rect -64 -102 -60 -98
rect -64 -110 -60 -106
rect -48 -106 -44 -102
rect -111 -118 -107 -114
rect -67 -118 -63 -114
rect -111 -126 -107 -122
rect -63 -126 -59 -122
rect -64 -134 -60 -130
rect -64 -142 -60 -138
rect -64 -150 -60 -146
rect -67 -158 -63 -154
rect -63 -166 -59 -162
rect -64 -174 -60 -170
rect -48 -178 -44 -174
rect -64 -182 -60 -178
rect -64 -190 -60 -186
rect -48 -186 -44 -182
<< m2contact >>
rect -73 18 -68 22
rect -73 -22 -68 -18
rect -119 -38 -115 -34
rect -73 -62 -68 -58
rect -119 -78 -115 -74
rect -73 -102 -68 -98
rect -119 -118 -115 -114
rect -73 -142 -68 -138
rect -119 -177 -115 -173
rect -73 -182 -68 -178
<< psubstratepcontact >>
rect -89 18 -85 22
rect -89 -22 -85 -18
rect -89 -62 -85 -58
rect -89 -102 -85 -98
rect -89 -142 -85 -138
rect -89 -182 -85 -178
<< nsubstratencontact >>
rect -56 18 -52 22
rect -56 -22 -52 -18
rect -56 -62 -52 -58
rect -56 -102 -52 -98
rect -56 -142 -52 -138
rect -56 -182 -52 -178
<< labels >>
rlabel metal1 -59 34 -57 37 1 Vdd
rlabel metal1 -88 42 -87 42 3 GND
rlabel metal1 -26 43 -24 44 7 GND
rlabel metal1 -18 45 -14 46 5 A
rlabel metal1 -11 45 -7 46 6 B
rlabel metal1 -59 -6 -57 -3 1 Vdd
rlabel metal1 -26 3 -24 4 7 GND
rlabel metal1 -18 5 -14 6 5 A
rlabel metal1 -11 5 -7 6 6 B
rlabel metal1 -59 -46 -57 -43 1 Vdd
rlabel metal1 -88 -38 -87 -38 3 GND
rlabel metal1 -26 -37 -24 -36 7 GND
rlabel metal1 -18 -35 -14 -34 5 A
rlabel metal1 -11 -35 -7 -34 6 B
rlabel metal1 -59 -86 -57 -83 1 Vdd
rlabel metal1 -88 -78 -87 -78 3 GND
rlabel metal1 -18 -75 -14 -74 5 A
rlabel metal1 -11 -75 -7 -74 6 B
rlabel metal1 -59 -126 -57 -123 1 Vdd
rlabel metal1 -88 -118 -87 -118 3 GND
rlabel metal1 -18 -115 -14 -114 5 A
rlabel metal1 -11 -115 -7 -114 6 B
rlabel metal1 -59 -166 -57 -163 1 Vdd
rlabel metal1 -88 -158 -87 -158 3 GND
rlabel metal1 -18 -155 -14 -154 5 A
rlabel metal1 -11 -155 -7 -154 6 B
rlabel metal1 -119 -190 -115 -188 2 Vdd
rlabel metal1 -120 -155 -120 -151 3 inbit
rlabel metal1 -120 -94 -120 -90 3 s0
rlabel metal1 -120 -54 -120 -50 3 s1
rlabel metal1 -120 45 -120 49 4 load
rlabel metal1 -120 -134 -120 -130 3 shift
rlabel metal1 -120 5 -120 9 3 add
<< end >>
