magic
tech scmos
timestamp 1428729551
<< pwell >>
rect -105 -16 -69 -1
rect -52 -16 -27 1
rect -103 -18 -73 -16
<< nwell >>
rect -100 16 -90 19
rect -100 15 -77 16
rect -100 5 -37 15
<< polysilicon >>
rect -58 25 -54 27
rect -92 23 -54 25
rect -92 12 -90 23
rect -50 18 -28 20
rect -50 14 -48 18
rect -42 14 -40 16
rect -84 12 -82 14
rect -110 5 -98 7
rect -110 4 -108 5
rect -100 -22 -98 5
rect -92 1 -90 8
rect -84 5 -82 8
rect -84 3 -74 5
rect -92 -1 -82 1
rect -92 -8 -90 -6
rect -84 -8 -82 -1
rect -76 -3 -74 3
rect -50 3 -48 10
rect -42 7 -40 10
rect -42 5 -20 7
rect -50 1 -40 3
rect -76 -5 -65 -3
rect -92 -15 -90 -12
rect -84 -14 -82 -12
rect -76 -16 -74 -5
rect -67 -12 -65 -5
rect -50 -6 -48 -4
rect -42 -6 -40 1
rect -67 -14 -60 -12
rect -50 -14 -48 -10
rect -42 -12 -40 -10
rect -34 -12 -32 5
rect -22 4 -20 5
rect -38 -14 -32 -12
rect -89 -18 -74 -16
rect -72 -22 -70 -19
rect -62 -21 -60 -14
rect -53 -16 -48 -14
rect -42 -16 -36 -14
rect -50 -18 -40 -16
rect -34 -19 -26 -17
rect -34 -20 -32 -19
rect -48 -21 -32 -20
rect -100 -24 -70 -22
rect -62 -22 -32 -21
rect -62 -23 -46 -22
<< ndiffusion >>
rect -93 -12 -92 -8
rect -90 -12 -89 -8
rect -85 -12 -84 -8
rect -82 -12 -81 -8
rect -51 -10 -50 -6
rect -48 -10 -47 -6
rect -43 -10 -42 -6
rect -40 -10 -39 -6
<< pdiffusion >>
rect -93 8 -92 12
rect -90 8 -89 12
rect -85 8 -84 12
rect -82 8 -81 12
rect -51 10 -50 14
rect -48 10 -47 14
rect -43 10 -42 14
rect -40 10 -39 14
<< metal1 >>
rect -140 27 -58 31
rect -54 27 64 31
rect -140 18 -28 22
rect -24 18 64 22
rect -101 8 -97 12
rect -77 8 -73 12
rect -59 10 -55 14
rect -35 10 -31 14
rect -47 9 -43 10
rect -89 7 -85 8
rect -140 0 -112 4
rect -77 -2 -63 2
rect -18 0 64 4
rect -47 -6 -43 -5
rect -89 -8 -85 -7
rect -101 -12 -97 -8
rect -77 -12 -73 -8
rect -59 -10 -55 -6
rect -35 -10 -31 -6
rect -47 -11 -43 -10
rect -140 -19 -93 -15
rect -66 -18 -57 -14
rect -66 -21 -62 -18
rect -22 -19 64 -15
<< metal2 >>
rect -82 27 -51 31
rect -105 12 -101 26
rect -82 22 -78 27
rect -82 18 -69 22
rect -105 -8 -101 8
rect -73 12 -69 18
rect -89 2 -85 3
rect -89 -2 -81 2
rect -89 -3 -85 -2
rect -89 -8 -85 -7
rect -73 -8 -69 8
rect -63 14 -59 15
rect -63 2 -59 10
rect -63 -6 -59 -2
rect -47 9 -43 10
rect -47 -1 -43 5
rect -47 -6 -43 -5
rect -31 -6 -27 10
rect -53 -15 -47 -14
rect -53 -18 -43 -15
rect -53 -19 -49 -18
rect -90 -23 -49 -19
rect -90 -27 -86 -23
<< ntransistor >>
rect -92 -12 -90 -8
rect -84 -12 -82 -8
rect -50 -10 -48 -6
rect -42 -10 -40 -6
<< ptransistor >>
rect -92 8 -90 12
rect -84 8 -82 12
rect -50 10 -48 14
rect -42 10 -40 14
<< polycontact >>
rect -58 27 -54 31
rect -28 18 -24 22
rect -112 0 -108 4
rect -93 -19 -89 -15
rect -22 0 -18 4
rect -70 -21 -66 -17
rect -57 -18 -53 -14
rect -26 -19 -22 -15
<< ndcontact >>
rect -97 -12 -93 -8
rect -89 -12 -85 -8
rect -81 -12 -77 -8
rect -55 -10 -51 -6
rect -47 -10 -43 -6
rect -39 -10 -35 -6
<< pdcontact >>
rect -97 8 -93 12
rect -89 8 -85 12
rect -81 8 -77 12
rect -55 10 -51 14
rect -47 10 -43 14
rect -39 10 -35 14
<< m2contact >>
rect -105 8 -101 12
rect -73 8 -69 12
rect -63 10 -59 14
rect -31 10 -27 14
rect -89 3 -85 7
rect -47 5 -43 9
rect -81 -2 -77 2
rect -63 -2 -59 2
rect -89 -7 -85 -3
rect -47 -5 -43 -1
rect -105 -12 -101 -8
rect -73 -12 -69 -8
rect -63 -10 -59 -6
rect -31 -10 -27 -6
rect -47 -15 -43 -11
<< psubstratepcontact >>
rect -105 -5 -101 -1
rect -31 -3 -27 1
<< end >>
