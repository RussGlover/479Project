magic
tech scmos
timestamp 1427503788
<< pwell >>
rect -85 33 -72 46
rect -89 9 -73 33
<< nwell >>
rect -68 9 -52 46
<< polysilicon >>
rect -91 48 -51 49
rect -91 47 -74 48
rect -70 47 -51 48
rect -83 39 -81 41
rect -77 39 -67 41
rect -59 39 -57 41
rect -72 33 -70 39
rect -90 23 -81 25
rect -77 23 -64 25
rect -60 23 -52 25
rect -90 15 -81 17
rect -77 15 -64 17
rect -60 15 -52 17
<< ndiffusion >>
rect -81 41 -77 42
rect -81 38 -77 39
rect -81 25 -77 26
rect -81 17 -77 23
rect -81 14 -77 15
rect -81 9 -77 10
<< pdiffusion >>
rect -63 42 -59 46
rect -67 41 -59 42
rect -67 38 -59 39
rect -67 34 -63 38
rect -64 25 -60 26
rect -64 22 -60 23
rect -64 17 -60 18
rect -64 14 -60 15
rect -64 9 -60 10
<< metal1 >>
rect -77 44 -74 46
rect -70 44 -67 46
rect -77 42 -67 44
rect -85 34 -81 38
rect -59 34 -56 38
rect -77 29 -73 30
rect -69 29 -68 33
rect -77 26 -68 29
rect -60 26 -56 30
rect -73 22 -68 26
rect -68 18 -64 22
rect -85 10 -81 14
rect -60 10 -56 14
<< metal2 >>
rect -89 38 -85 46
rect -89 14 -85 34
rect -56 38 -52 46
rect -56 30 -52 34
rect -89 9 -85 10
rect -56 14 -52 26
rect -56 9 -52 10
<< ntransistor >>
rect -81 39 -77 41
rect -81 23 -77 25
rect -81 15 -77 17
<< ptransistor >>
rect -67 39 -59 41
rect -64 23 -60 25
rect -64 15 -60 17
<< polycontact >>
rect -74 44 -70 48
rect -73 29 -69 33
<< ndcontact >>
rect -81 42 -77 46
rect -81 34 -77 38
rect -81 26 -77 30
rect -81 10 -77 14
<< pdcontact >>
rect -67 42 -63 46
rect -63 34 -59 38
rect -64 26 -60 30
rect -64 18 -60 22
rect -64 10 -60 14
<< m2contact >>
rect -89 34 -85 38
rect -56 34 -52 38
rect -56 26 -52 30
rect -73 18 -68 22
rect -89 10 -85 14
rect -56 10 -52 14
<< psubstratepcontact >>
rect -89 18 -85 22
<< nsubstratencontact >>
rect -56 18 -52 22
<< labels >>
rlabel polysilicon -90 23 -81 25 3 A
rlabel polysilicon -90 15 -81 17 3 B
rlabel metal2 -89 14 -85 37 3 GND
rlabel polysilicon -91 47 -51 49 5 out
rlabel metal2 -56 38 -52 46 7 Vdd
<< end >>
