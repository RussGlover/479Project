magic
tech scmos
timestamp 1428965811
<< pwell >>
rect 554 -143 570 193
rect 1003 162 1069 175
rect 1003 130 1019 162
<< nwell >>
rect 575 -142 591 177
rect 1024 135 1068 160
<< polysilicon >>
rect 546 193 552 195
rect 549 139 551 193
rect 601 171 603 177
rect 591 169 603 171
rect 1033 170 1035 232
rect 1057 170 1059 220
rect 587 161 599 163
rect 597 147 599 161
rect 1033 156 1035 166
rect 1057 156 1059 166
rect 1033 150 1035 152
rect 1057 150 1059 152
rect 597 145 617 147
rect 549 137 562 139
rect 566 137 579 139
rect 583 137 585 139
rect 560 113 562 115
rect 566 113 579 115
rect 583 113 605 115
rect 560 -49 562 -47
rect 566 -49 579 -47
rect 583 -49 595 -47
rect 560 -66 562 -64
rect 566 -66 579 -64
rect 583 -66 603 -64
rect 612 -131 614 -107
rect 560 -133 562 -131
rect 566 -133 579 -131
rect 583 -133 614 -131
<< ndiffusion >>
rect 1032 166 1033 170
rect 1035 166 1036 170
rect 1056 166 1057 170
rect 1059 166 1060 170
rect 562 139 566 140
rect 562 136 566 137
rect 562 115 566 116
rect 562 112 566 113
rect 562 -47 566 -46
rect 562 -50 566 -49
rect 562 -64 566 -63
rect 562 -67 566 -66
rect 562 -131 566 -130
rect 562 -134 566 -133
<< pdiffusion >>
rect 1032 152 1033 156
rect 1035 152 1036 156
rect 1056 152 1057 156
rect 1059 152 1060 156
rect 579 139 583 140
rect 579 136 583 137
rect 579 115 583 116
rect 579 112 583 113
rect 579 -47 583 -46
rect 579 -50 583 -49
rect 579 -64 583 -63
rect 579 -67 583 -66
rect 579 -131 583 -130
rect 579 -134 583 -133
<< metal1 >>
rect -2554 246 599 250
rect 595 228 599 246
rect 633 240 690 244
rect 625 232 1032 236
rect 595 224 1092 228
rect 533 217 605 221
rect 533 210 816 214
rect 535 203 613 207
rect 617 203 824 207
rect 503 191 542 195
rect 604 177 605 181
rect 999 174 1056 178
rect 1028 170 1032 174
rect 1052 170 1056 174
rect 609 161 808 165
rect 1036 163 1040 166
rect 1060 163 1064 166
rect 1036 159 1048 163
rect 690 157 767 158
rect 657 149 661 153
rect 694 154 767 157
rect 1036 156 1040 159
rect 690 148 694 153
rect 621 144 625 148
rect 511 140 562 144
rect 566 140 579 144
rect 558 132 562 136
rect 583 132 587 136
rect 763 130 767 154
rect 1028 148 1032 152
rect 970 144 1036 148
rect 970 134 974 144
rect 1036 139 1040 144
rect 914 130 974 134
rect 527 116 562 120
rect 566 116 579 120
rect 605 116 609 117
rect 558 108 562 112
rect 583 108 587 112
rect 607 104 625 108
rect 936 104 958 108
rect 936 84 940 104
rect 970 87 974 130
rect 1044 129 1048 159
rect 1060 159 1072 163
rect 1060 156 1064 159
rect 1052 148 1056 152
rect 1068 134 1072 159
rect 983 104 1004 108
rect 534 77 614 81
rect 531 55 603 59
rect 531 10 535 55
rect 603 45 622 49
rect 603 17 607 45
rect 917 28 937 32
rect 595 5 623 9
rect 558 -46 562 -42
rect 583 -46 587 -42
rect 595 -46 599 5
rect 535 -54 562 -50
rect 566 -54 579 -50
rect 595 -54 599 -50
rect 535 -63 562 -59
rect 566 -63 579 -59
rect 603 -63 607 -3
rect 558 -71 562 -67
rect 583 -71 587 -67
rect 603 -77 607 -67
rect 530 -81 607 -77
rect 611 -35 622 -31
rect 531 -89 595 -85
rect 531 -100 535 -89
rect 611 -103 615 -35
rect 757 -38 761 -31
rect 548 -107 611 -103
rect 619 -56 625 -52
rect 619 -115 623 -56
rect 535 -119 623 -115
rect 558 -130 562 -126
rect 583 -130 587 -126
rect 535 -138 562 -134
rect 566 -138 579 -134
rect 535 -145 544 -141
rect 627 -148 631 -90
rect 657 -129 661 -91
rect 690 -148 694 -89
rect 720 -129 724 -90
rect 535 -152 694 -148
<< metal2 >>
rect -2331 246 -2327 254
rect -2118 246 -2114 254
rect -1905 246 -1901 254
rect -1692 246 -1688 254
rect -1479 246 -1475 254
rect -1266 246 -1262 254
rect -1053 246 -1049 254
rect -831 246 -827 254
rect -658 246 -654 254
rect -484 246 -480 254
rect -310 246 -306 254
rect -137 246 -133 254
rect 37 246 41 254
rect 212 246 216 254
rect 386 246 390 254
rect -2558 39 -2554 246
rect -2558 35 -2553 39
rect -2201 -156 -2197 -132
rect -1988 -156 -1984 -132
rect -1775 -156 -1771 -132
rect -1562 -156 -1558 -132
rect -1349 -156 -1345 -132
rect -1136 -156 -1132 -132
rect -923 -156 -919 -132
rect -734 -156 -730 -37
rect -561 -156 -557 -37
rect -387 -155 -383 -34
rect -213 -156 -209 -39
rect -40 -156 -36 -39
rect 134 -156 138 -40
rect 309 -156 313 -40
rect 483 -156 487 -36
rect 491 -42 495 239
rect 499 195 503 231
rect 507 144 511 224
rect 605 221 609 254
rect 523 120 527 210
rect 605 181 609 217
rect 613 207 617 254
rect 621 236 625 254
rect 629 244 633 254
rect 637 221 641 254
rect 641 217 661 221
rect 605 165 609 177
rect 554 136 558 151
rect 554 112 558 132
rect 491 -148 495 -46
rect 501 -108 505 77
rect 554 -42 558 108
rect 554 -67 558 -46
rect 544 -141 548 -107
rect 554 -126 558 -71
rect 587 136 591 151
rect 587 112 591 132
rect 605 121 609 161
rect 657 157 661 217
rect 690 157 694 240
rect 808 112 812 161
rect 587 -42 591 108
rect 603 59 607 104
rect 816 105 820 210
rect 824 98 828 203
rect 995 127 999 174
rect 1040 144 1052 148
rect 1092 141 1096 224
rect 995 123 1003 127
rect 962 104 979 108
rect 603 1 607 13
rect 587 -67 591 -46
rect 587 -126 591 -71
rect 595 -85 599 -58
rect 614 -129 618 77
rect 704 -42 757 -38
rect 704 -129 708 -42
rect 614 -133 657 -129
rect 661 -133 720 -129
<< ntransistor >>
rect 1033 166 1035 170
rect 1057 166 1059 170
rect 562 137 566 139
rect 562 113 566 115
rect 562 -49 566 -47
rect 562 -66 566 -64
rect 562 -133 566 -131
<< ptransistor >>
rect 1033 152 1035 156
rect 1057 152 1059 156
rect 579 137 583 139
rect 579 113 583 115
rect 579 -49 583 -47
rect 579 -66 583 -64
rect 579 -133 583 -131
<< polycontact >>
rect 1032 232 1036 236
rect 542 191 546 195
rect 600 177 604 181
rect 1056 220 1060 224
rect 617 144 621 148
rect 605 112 609 116
rect 595 -50 599 -46
rect 603 -67 607 -63
rect 611 -107 615 -103
<< ndcontact >>
rect 1028 166 1032 170
rect 1036 166 1040 170
rect 1052 166 1056 170
rect 1060 166 1064 170
rect 562 140 566 144
rect 562 132 566 136
rect 562 116 566 120
rect 562 108 566 112
rect 562 -46 566 -42
rect 562 -54 566 -50
rect 562 -63 566 -59
rect 562 -71 566 -67
rect 562 -130 566 -126
rect 562 -138 566 -134
<< pdcontact >>
rect 1028 152 1032 156
rect 1036 152 1040 156
rect 1052 152 1056 156
rect 1060 152 1064 156
rect 579 140 583 144
rect 579 132 583 136
rect 579 116 583 120
rect 579 108 583 112
rect 579 -46 583 -42
rect 579 -54 583 -50
rect 579 -63 583 -59
rect 579 -71 583 -67
rect 579 -130 583 -126
rect 579 -138 583 -134
<< m2contact >>
rect -2558 246 -2554 250
rect 491 239 495 243
rect 499 231 503 235
rect 629 240 633 244
rect 690 240 694 244
rect 621 232 625 236
rect 507 224 511 228
rect 1092 224 1096 228
rect 605 217 609 221
rect 637 217 641 221
rect 523 210 527 214
rect 816 210 820 214
rect 613 203 617 207
rect 824 203 828 207
rect 499 191 503 195
rect 605 177 609 181
rect 995 174 999 178
rect 605 161 609 165
rect 808 161 812 165
rect 554 151 558 155
rect 587 151 591 155
rect 657 153 661 157
rect 690 153 694 157
rect 507 140 511 144
rect 554 132 558 136
rect 587 132 591 136
rect 1036 144 1040 148
rect 523 116 527 120
rect 605 117 609 121
rect 554 108 558 112
rect 587 108 591 112
rect 808 108 812 112
rect 603 104 607 108
rect 816 101 820 105
rect 958 104 962 108
rect 824 94 828 98
rect 1052 144 1056 148
rect 1092 137 1096 141
rect 1003 123 1007 127
rect 979 104 983 108
rect 501 77 505 81
rect 614 77 618 81
rect 603 55 607 59
rect 603 13 607 17
rect 491 -46 495 -42
rect 554 -46 558 -42
rect 587 -46 591 -42
rect 595 -58 599 -54
rect 603 -3 607 1
rect 554 -71 558 -67
rect 587 -71 591 -67
rect 595 -89 599 -85
rect 987 -34 991 -30
rect 757 -42 761 -38
rect 544 -107 548 -103
rect 501 -112 505 -108
rect 994 -86 998 -82
rect 554 -130 558 -126
rect 587 -130 591 -126
rect 544 -145 548 -141
rect 657 -133 661 -129
rect 720 -133 724 -129
rect 491 -152 495 -148
use dp8  dp8_0
timestamp 1428827926
transform 1 0 -1088 0 1 -152
box -1491 0 1623 399
use andgate  andgate_0
timestamp 1428729313
transform 1 0 648 0 1 146
box -96 9 -57 49
use inputCombLogic2  inputCombLogic2_0
timestamp 1428802844
transform 1 0 1077 0 1 -184
box -455 90 19 333
<< labels >>
rlabel metal2 -2331 253 -2327 254 5 divisorin_6
rlabel metal2 -2118 253 -2114 254 5 divisorin_5
rlabel metal2 -1905 253 -1901 254 5 divisorin_4
rlabel metal2 -1479 253 -1475 254 5 divisorin_2
rlabel metal2 -1053 253 -1049 254 5 divisorin_0
rlabel metal2 -1266 253 -1262 254 5 divisorin_1
rlabel metal2 -1692 253 -1688 254 5 divisorin_3
rlabel metal2 -831 253 -827 254 5 dividendin_7
rlabel metal2 -658 253 -654 254 5 dividendin_6
rlabel metal2 -484 253 -480 254 5 dividendin_5
rlabel metal2 -310 253 -306 254 5 dividendin_4
rlabel metal2 -137 253 -133 254 5 dividendin_3
rlabel metal2 37 253 41 254 5 dividendin_2
rlabel metal2 212 253 216 254 5 dividendin_1
rlabel metal2 386 253 390 254 5 dividendin_0
rlabel metal2 -2201 -156 -2197 -155 1 remainder_6
rlabel metal2 -1988 -156 -1984 -155 1 remainder_5
rlabel metal2 -1775 -156 -1771 -155 1 remainder_4
rlabel metal2 -1562 -156 -1558 -155 1 remainder_3
rlabel metal2 -1349 -156 -1345 -155 1 remainder_2
rlabel metal2 -1136 -156 -1132 -155 1 remainder_1
rlabel metal2 -923 -156 -919 -155 1 remainder_0
rlabel metal2 -734 -156 -730 -155 1 quotient_7
rlabel metal2 -561 -156 -557 -155 1 quotient_6
rlabel metal2 -387 -155 -383 -154 1 quotient_5
rlabel metal2 -213 -156 -209 -155 1 quotient_4
rlabel metal2 -40 -156 -36 -155 1 quotient_3
rlabel metal2 134 -156 138 -155 1 quotient_2
rlabel metal2 309 -156 313 -155 1 quotient_1
rlabel metal2 483 -156 487 -155 1 quotient_0
rlabel metal2 629 253 633 254 5 Vdd
rlabel metal2 613 253 617 254 5 reset
rlabel metal2 605 253 609 254 5 clk
rlabel metal2 621 253 625 254 5 start
rlabel metal2 637 253 641 254 5 GND
<< end >>
